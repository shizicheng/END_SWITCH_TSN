module dmac_mng #(
        parameter                           PORT_NUM                =      8                                    ,   // �������Ķ˿�??
        parameter                           HASH_DATA_WIDTH         =      15                                   ,   // ��ϣ�����???��λ��֧??32K??
        parameter                           REG_ADDR_BUS_WIDTH      =      8                                    ,   // ���� MAC ������üĴ�����??λ��
        parameter                           REG_DATA_BUS_WIDTH      =      16                                   ,   // ���� MAC ������üĴ�������λ??
        parameter                           PORT_NUM_BIT            =      clog2(PORT_NUM)                      ,   // �˿ں�λ??
        parameter                           MAC_TABLE_DEPTH         =      2**HASH_DATA_WIDTH                   ,   // MAC����ȣ�32K
        parameter                           AGE_TIME_WIDTH          =      10                                   ,   // �ϻ�ʱ��λ��֧??1024??
        parameter                           VLAN_ID_WIDTH           =      12                                   ,   // VLAN IDλ��
        parameter                           MAC_ADDR_WIDTH          =      48                                   ,   // MAC��ַλ��
        parameter                           CLK_FREQ_MHZ            =      250                                  ,   // ����ʱ��Ƶ�� 
        parameter                           TABLE_FULL_THRESHOLD    =      29491                                ,   // MAC������???��90% of 32K = 29491??
        parameter                           ENTRY_WIDTH             =      1 + AGE_TIME_WIDTH + VLAN_ID_WIDTH 
                                                                           + PORT_NUM + MAC_ADDR_WIDTH          ,   // ����λ��: [��Чλ[1] + �ϻ�ʱ��[AGE_TIME_WIDTH-1:0] + VLAN_ID[VLAN_ID_WIDTH-1:0] + �˿ں�[PORT_NUM-1:0] + MAC��ַ[MAC_ADDR_WIDTH-1:0]]
        parameter                           AGE_SCAN_INTERVAL       =      5                                    ,   // �ϻ�ɨ��������??
        parameter                           SIM_MODE                =      0                                        // ����ģʽ??1=��???����ģʽ��0=����ģʽ
)(                      
        input               wire                                        i_clk                                   ,
        input               wire                                        i_rst                                   , 
        /*----------------------------- �Ĵ���д���ƽӿ� ------------------------------*/     
        //input               wire                                        i_reg_bus_we                            , // �Ĵ���дʹ��
        //input               wire        [REG_ADDR_BUS_WIDTH-1:0]        i_reg_bus_addr                          , // �Ĵ���д��ַ
        //input               wire        [REG_DATA_BUS_WIDTH-1:0]        i_reg_bus_data                          , // �Ĵ���д����
        //input               wire                                        i_reg_bus_data_vld                      , // �Ĵ���д����ʹ��
        
        /*----------------------------- �Ĵ��������ƽӿ� ------------------------------*/
        //input               wire                                        i_reg_bus_re                            , // �Ĵ�����ʹ��
        //input               wire        [REG_ADDR_BUS_WIDTH-1:0]        i_reg_bus_raddr                         , // �Ĵ�������ַ
        //output              wire        [REG_DATA_BUS_WIDTH-1:0]        o_reg_bus_rdata                         , // �Ĵ���������
        //output              wire                                        o_reg_bus_rdata_vld                     , // �Ĵ�����������Ч
        
        /*----------------------------- DMAC/SMAC ���ӿ� ------------------------------*/
        input               wire        [VLAN_ID_WIDTH-1:0]             i_vlan_id                               , // ���뱨�ĵ�VLAN ID
        input               wire        [MAC_ADDR_WIDTH-1:0]            i_dmac                                  , // Ŀ��MAC��ַ����
        input               wire        [HASH_DATA_WIDTH-1:0]           i_dmac_hash_addr                        , // Ŀ��MAC��hash��ַ
        input               wire                                        i_dmac_hash_vld                         , // DMAC hash��������Ч  
        input               wire        [MAC_ADDR_WIDTH-1:0]            i_smac                                  , // ԴMAC��ַ����
        input               wire        [HASH_DATA_WIDTH-1:0]           i_smac_hash_addr                        , // ԴMAC��hash��ַ
        input               wire                                        i_smac_hash_vld                         , // SMAC hash��������Ч  
        input               wire        [PORT_NUM-1:0]                  i_rx_port                               , // ���ն˿�bitmap,ÿ��bit����??����??
        
        /*----------------------------- �������ӿ� ------------------------------*/                           
        output              wire                                        o_dmac_lookup_vld                       , // DMAC�������Ч
        output              wire        [PORT_NUM-1:0]                  o_dmac_tx_port                          , // DMAC�������ת����?? 
        output              wire                                        o_dmac_lookup_hit                       , // DMAC������б�־
        output              wire                                        o_lookup_clash                          , // ����ͻ��־����ϣ��??�б��MAC/VLAN��ƥ??
        output              wire                                        o_table_full                            , // MAC������־

        output              wire        [HASH_DATA_WIDTH-1:0]           o_mac_table_addr                        ,
        output              wire        [3:0]                           o_fsm_cur_state                         ,

        input               wire                                        i_table_clear_req                       ,
        input               wire        [AGE_TIME_WIDTH-1:0]            i_age_time_threshold                    ,
        input               wire                                        i_table_rd                              ,
        input               wire        [11:0]                          i_table_raddr                           ,
        input              wire         [14:0]                          i_table_full_threshold                  ,
        input              wire         [31:0]                          i_age_scan_interval                     , // �ϻ�ɨ�������üĴ������룩

        output              wire        [57:0]                          o_dmac_list_dout                        ,
        output              wire        [15:0]                          o_dmac_list_cnt                         ,
        output              wire                                        o_dmac_list_full_er_stat                ,
        output              wire        [15:0]                          o_dmac_list_full_er_cnt                 ,

        output              wire        [14:0]                          o_table_entry_cnt                       ,
        output              wire        [15:0]                          o_learn_success_cnt                     ,
        output              wire        [REG_DATA_BUS_WIDTH-1:0]        o_collision_cnt                         ,
        output              wire        [REG_DATA_BUS_WIDTH-1:0]        o_port_move_cnt                        
);

/*---------------------------------------- clog2���㺯�� -------------------------------------------*/
function integer clog2;
    input integer value;
    integer temp;
    begin
        temp = value - 1;
        for (clog2 = 0; temp > 0; clog2 = clog2 + 1)
            temp = temp >> 1;
    end
endfunction 

/*---------------------------------------- �Ĵ�����??���� -------------------------------------------*/
//localparam  REG_AGE_TIME_THRESHOLD      = 8'h00                             ; // �ϻ�ʱ����???���üĴ���
//localparam  REG_TABLE_CLEAR             = 8'h01                             ; // MAC����ռĴ���
//localparam  REG_TABLE_FULL_THRESHOLD    = 8'h02                             ; // MAC������???���üĴ���
//localparam  REG_AGE_SCAN_INTERVAL       = 8'h03                             ; // �ϻ�ɨ�������üĴ�??
//localparam  REG_TABLE_ENTRY_cnt         = 8'h04                             ; // MAC�����������ֻ��??
//localparam  REG_LEARN_STATISTICS        = 8'h05                             ; // MACѧϰͳ�ƼĴ�����ֻ��??
//localparam  REG_COLLISION_STATISTICS    = 8'h06                             ; // ��ϣ��ͻͳ�ƼĴ�����ֻ��??
//localparam  REG_PORT_MOVE_STATISTICS    = 8'h07                             ; // �˿��ƶ�ͳ�ƼĴ�����ֻ��??

/*---------------------------------------- ״???������ -------------------------------------------*/
localparam  IDLE                        = 4'd0                              ; // ����״???
localparam  FIFO_READ_WAIT              = 4'd1                              ; // FIFO��ȡ�ȴ�״???��STDģʽ??Ҫ��
localparam  DMAC_LOOKUP                 = 4'd2                              ; // DMAC���״???
localparam  DMAC_REFRESH                = 4'd3                              ; // DMAC�����ϻ�ʱ��ˢ��״???
localparam  SMAC_LEARN_CHECK            = 4'd4                              ; // SMACѧϰ??��״??
localparam  SMAC_LEARN_UPDATE           = 4'd5                              ; // SMACѧϰ����״???
localparam  AGE_SCAN                    = 4'd6                              ; // �ϻ�ɨ��״???
localparam  AGE_UPDATE                  = 4'd7                              ; // �ϻ�����״???

/*---------------------------------------- �ڲ��źŶ��� -------------------------------------------*/
// ��������FIFO��ز�������??
localparam  INPUT_FIFO_DEPTH            = 8                                 ; // ����FIFO��ȣ�֧??8�����Ļ�??
localparam  INPUT_DATA_WIDTH            = VLAN_ID_WIDTH + MAC_ADDR_WIDTH*2 + 
                                          HASH_DATA_WIDTH*2 + 2 + PORT_NUM_BIT ; // ��������λ��VLAN+DMAC+SMAC+DMAC_HASH+SMAC_HASH+2��VLD+PORT

// 5������FIFO��λ��??
localparam  FIFO1_WIDTH                 = VLAN_ID_WIDTH + PORT_NUM         ; // FIFO1: VLAN_ID + RX_PORT(bitmap)
localparam  FIFO2_WIDTH                 = MAC_ADDR_WIDTH                    ; // FIFO2: DMAC
localparam  FIFO3_WIDTH                 = MAC_ADDR_WIDTH                    ; // FIFO3: SMAC  
localparam  FIFO4_WIDTH                 = HASH_DATA_WIDTH + 1               ; // FIFO4: DMAC_HASH_ADDR + DMAC_HASH_VLD
localparam  FIFO5_WIDTH                 = HASH_DATA_WIDTH + 1               ; // FIFO5: SMAC_HASH_ADDR + SMAC_HASH_VLD

// 5������FIFO�Ľӿ���??
// FIFO1: VLAN_ID + RX_PORT
wire                                    w_fifo1_wr_en                       ; // FIFO1дʹ??
wire        [FIFO1_WIDTH-1:0]           w_fifo1_din                         ; // FIFO1��������
wire                                    w_fifo1_full                        ; // FIFO1����??
wire                                    w_fifo1_rd_en                       ; // FIFO1��ʹ??
wire        [FIFO1_WIDTH-1:0]           w_fifo1_dout                        ; // FIFO1�������
wire                                    w_fifo1_empty                       ; // FIFO1�ձ�??

// FIFO2: DMAC
wire                                    w_fifo2_wr_en                       ; // FIFO2дʹ??
wire        [FIFO2_WIDTH-1:0]           w_fifo2_din                         ; // FIFO2��������
wire                                    w_fifo2_full                        ; // FIFO2����??
wire                                    w_fifo2_rd_en                       ; // FIFO2��ʹ??
wire        [FIFO2_WIDTH-1:0]           w_fifo2_dout                        ; // FIFO2�������
wire                                    w_fifo2_empty                       ; // FIFO2�ձ�??

// FIFO3: SMAC  
wire                                    w_fifo3_wr_en                       ; // FIFO3дʹ??
wire        [FIFO3_WIDTH-1:0]           w_fifo3_din                         ; // FIFO3��������
wire                                    w_fifo3_full                        ; // FIFO3����??
wire                                    w_fifo3_rd_en                       ; // FIFO3��ʹ??
wire        [FIFO3_WIDTH-1:0]           w_fifo3_dout                        ; // FIFO3�������
wire                                    w_fifo3_empty                       ; // FIFO3�ձ�??

// FIFO4: DMAC_HASH_ADDR + DMAC_HASH_VLD
wire                                    w_fifo4_wr_en                       ; // FIFO4дʹ??
wire        [FIFO4_WIDTH-1:0]           w_fifo4_din                         ; // FIFO4��������
wire                                    w_fifo4_full                        ; // FIFO4����??
wire                                    w_fifo4_rd_en                       ; // FIFO4��ʹ??
wire        [FIFO4_WIDTH-1:0]           w_fifo4_dout                        ; // FIFO4�������
wire                                    w_fifo4_empty                       ; // FIFO4�ձ�??

// FIFO5: SMAC_HASH_ADDR + SMAC_HASH_VLD
wire                                    w_fifo5_wr_en                       ; // FIFO5дʹ??
wire        [FIFO5_WIDTH-1:0]           w_fifo5_din                         ; // FIFO5��������
wire                                    w_fifo5_full                        ; // FIFO5����??
wire                                    w_fifo5_rd_en                       ; // FIFO5��ʹ??
wire        [FIFO5_WIDTH-1:0]           w_fifo5_dout                        ; // FIFO5�������
wire                                    w_fifo5_empty                       ; // FIFO5�ձ�??

// �ۺ�FIFO״???��??
wire                                    w_all_fifo_full                     ; // ??��FIFO����??
wire                                    w_all_fifo_empty                    ; // ??��FIFO�ձ�??

// ��FIFO��������н���������??
wire        [VLAN_ID_WIDTH-1:0]         w_fifo_vlan_id                      ;
wire        [MAC_ADDR_WIDTH-1:0]        w_fifo_dmac                         ;
wire        [MAC_ADDR_WIDTH-1:0]        w_fifo_smac                         ;
wire        [HASH_DATA_WIDTH-1:0]       w_fifo_dmac_hash_addr               ;       
wire        [HASH_DATA_WIDTH-1:0]       w_fifo_smac_hash_addr               ;
wire        [PORT_NUM-1:0]              w_fifo_rx_port                      ; // ���ն˿�bitmap

// �Ĵ��������??  
//reg                                     r_reg_bus_we                        ;
//reg         [REG_ADDR_BUS_WIDTH-1:0]    r_reg_bus_addr                      ;
//reg         [REG_DATA_BUS_WIDTH-1:0]    r_reg_bus_data                      ;
//reg                                     r_reg_bus_data_vld                  ;

// �Ĵ����������ź�
//reg                                     r_reg_bus_re                        ;
//reg         [REG_ADDR_BUS_WIDTH-1:0]    r_reg_bus_raddr                     ;
//reg         [REG_DATA_BUS_WIDTH-1:0]    r_reg_bus_rdata                     ;
//reg                                     r_reg_bus_rdata_vld                 ;

// ����Ĵ�??
reg                                     r_dmac_lookup_vld                   ;
reg         [PORT_NUM-1:0]              r_dmac_tx_port                      ;             
reg                                     r_dmac_lookup_hit                   ;
reg                                     r_lookup_clash                      ; // ����ͻ��־�Ĵ�??

// ״???�����
reg         [3:0]                       r_fsm_cur_state                     ;
reg         [3:0]                       r_fsm_nxt_state                     ;
reg         [15:0]                      r_state_cnt                         ; // ״???������������ÿ��״̬����ʱ??

// MAC��洢���ӿ�
reg         [HASH_DATA_WIDTH-1:0]       r_mac_table_addr                    ;
reg         [ENTRY_WIDTH-1:0]           r_mac_table_wdata                   ;
wire        [ENTRY_WIDTH-1:0]           w_mac_table_rdata                   ;
reg                                     r_mac_table_we                      ;
reg                                     r_mac_table_re                      ;

// �Ĵ�����ȡMAC��Ķ���ͨ��
reg         [HASH_DATA_WIDTH-1:0]       r_reg_table_raddr                   ; // �Ĵ��������??
reg                                     r_reg_table_rd                      ; // �Ĵ�������ʹ??


// ���üĴ�??
//reg         [AGE_TIME_WIDTH-1:0]        r_age_time_threshold                ; // �ϻ�ʱ����???��Ĭ��300�룩
//reg                                     r_table_clear_req                   ; // �������??
//reg         [14:0]                      r_table_full_threshold              ; // MAC������???���üĴ���
//reg         [31:0]                      r_age_scan_interval                 ; // �ϻ�ɨ�������üĴ������룩
reg                                       r_dmac_list_full_er_stat            ; // DMAC�б�������־
reg           [15:0]                      r_dmac_list_full_er_cnt             ; // DMAC�б���������??

// ͳ�ƼĴ�??
reg         [31:0]                      r_learn_success_cnt               ; // ѧϰ�ɹ�����??
reg         [31:0]                      r_learn_fail_cnt                  ; // ѧϰʧ�ܼ���??
reg         [31:0]                      r_collision_cnt                   ; // ��ϣ��ͻ����??
reg         [31:0]                      r_port_move_cnt                   ; // �˿��ƶ�����??

// ����������
reg         [14:0]                      r_table_entry_cnt                   ; // MAC����Ч�������������??32768??
reg                                     r_entry_add                         ; // ������ӱ�־
reg                                     r_entry_del                         ; // ����ɾ����־
wire                                    w_table_full                        ; // ����״???��??
wire                                    w_age_scan_trigger                  ; // �ϻ�ɨ�败���ź�
reg                                     r_table_full                        ; // ����״???��??
// �ϻ�����ź�
reg                                     r_age_scan_en                       ; // �ϻ�ɨ��ʹ��
reg                                     r_age_timer_pulse                   ; // �ϻ���ʱ�����壨1�����壩
reg         [AGE_TIME_WIDTH-1:0]        r_global_timestamp                  ; // ȫ��ʱ�������������??
reg         [7:0]                       r_clear_burst_cnt                   ; // ���ͻ������������������������??
reg                                     r_agescan_cnt                       ; // �ϻ���ַ���ּ���??
reg         [HASH_DATA_WIDTH-1:0]       r_age_scan_breakpoint               ; // �ϻ�ɨ��ϵ��ַ

// �ּ�ʱ������������??
reg         [15:0]                      r_us_cnt                            ; // ΢���������1-65535us��֧�ֲ�ͬʱ��Ƶ�ʣ�
reg         [9:0]                       r_ms_cnt                            ; // �������??
reg         [31:0]                      r_s_cnt                             ; // �����ܼ�������������??1���������ɣ�
reg         [31:0]                      r_age_scan_timer                    ; // �ϻ�ɨ�������������룩
reg                                     r_us_pulse                          ;  
reg                                     r_ms_pulse                          ;  

reg                                     r_can_use_direct_path               ;

// ʱ����� - ֧�ַ���ģʽ������ģ??
localparam  US_CNT_MAX                  = SIM_MODE ? 16'd5 : CLK_FREQ_MHZ   ; // ����ģʽ??10��ʱ����??=1us������ģʽ��CLK_FREQ_MHZ��ʱ����??=1us
localparam  MS_CNT_MAX                  = SIM_MODE ? 10'd5 : 10'd1000       ; // ����ģʽ??10us=1ms������ģʽ��1000us=1ms  
localparam  S_CNT_MAX                   = SIM_MODE ? 10'd5 : 10'd1000       ; // ����ģʽ??10ms=1s������ģʽ��1000ms=1s  
localparam  CLEAR_BURST_LIMIT           = 8'd16                             ; // ���ͻ�����ƣ�������??16����??����λ�����ݰ���??  

// ��������ź�
wire                                    w_entry_valid                       ; // ������Ч��־
wire        [AGE_TIME_WIDTH-1:0]        w_entry_age_time                    ; // �����ϻ�ʱ��
wire        [VLAN_ID_WIDTH-1:0]         w_entry_vlan_id                     ; // ����VLAN ID
wire        [PORT_NUM-1:0]              w_entry_port                        ; // ����˿ںţ�one-hot����??
wire        [MAC_ADDR_WIDTH-1:0]        w_entry_mac                         ; // ����MAC��ַ

// ���ƥ���ź�
wire                                    w_dmac_match                        ; // DMACƥ��
wire                                    w_smac_match                        ; // SMACƥ��
wire                                    w_smac_port_match                   ; // SMAC�˿�ƥ��
wire                                    w_entry_expired                     ; // ������ڱ�־

/*---------------------------------------- ��������FIFO���� -------------------------------------------*/
// �����ؼ��Ĵ���
reg                                     r_dmac_hash_vld_d1                  ; // DMAC��ϣ��Ч�ź��ӳ�????
reg                                     r_smac_hash_vld_d1                  ; // SMAC��ϣ��Ч�ź��ӳ�????
reg                                     r_entry_expired_flag                ;
// �����ؼ��???��
wire                                    w_dmac_hash_vld_posedge             ; // DMAC��ϣ��Ч����??
wire                                    w_smac_hash_vld_posedge             ; // SMAC��ϣ��Ч����??
wire                                    w_both_hash_valid                   ; // ����hash����??
wire                                    w_new_packet_arrival                ; // �±��ĵ�����??
wire                                    w_can_use_direct_path               ; // ����ʹ��ֱ��·���ź�
wire                                    w_fifo_dmac_hash_vld                ;
wire                                    w_fifo_smac_hash_vld                ;

assign w_dmac_hash_vld_posedge = i_dmac_hash_vld == 1'd1 && r_dmac_hash_vld_d1 == 1'd0 ? 1'd1 : 1'd0      ;
assign w_smac_hash_vld_posedge = i_smac_hash_vld == 1'd1 && r_smac_hash_vld_d1 == 1'd0 ? 1'd1 : 1'd0      ;
assign w_both_hash_valid = w_dmac_hash_vld_posedge == 1'd1 && w_smac_hash_vld_posedge == 1'd1 ? 1'd1 : 1'd0;
assign w_new_packet_arrival = w_both_hash_valid;

// �ۺ�FIFO״???��??
assign w_all_fifo_full =  (w_fifo1_full == 1'd1) || (w_fifo2_full == 1'd1) || (w_fifo3_full == 1'd1) || (w_fifo4_full == 1'd1) || (w_fifo5_full == 1'd1);
assign w_all_fifo_empty = (w_fifo1_empty == 1'd1) && (w_fifo2_empty == 1'd1) && (w_fifo3_empty == 1'd1) && (w_fifo4_empty == 1'd1) && (w_fifo5_empty == 1'd1);

// ֱ��·���жϣ�FIFOΪ����ģ�����ʱ����ֱ�Ӵ���
assign w_can_use_direct_path = w_new_packet_arrival == 1'd1 && w_all_fifo_empty == 1'd1 && i_table_clear_req == 1'd0 && r_fsm_cur_state == IDLE ? 1'd1 : 1'd0;

assign o_mac_table_addr                        = r_mac_table_addr;
assign o_fsm_cur_state                         = r_fsm_cur_state;
assign o_table_entry_cnt                       = r_table_entry_cnt;
assign o_learn_success_cnt                     = r_learn_success_cnt;
assign o_collision_cnt                         = r_collision_cnt;
assign o_port_move_cnt                         = r_port_move_cnt;  
assign o_dmac_list_full_er_cnt                 = r_dmac_list_full_er_cnt;
assign o_dmac_list_full_er_stat                = r_dmac_list_full_er_stat;
assign o_dmac_list_cnt                         = r_table_entry_cnt;




always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_dmac_hash_vld_d1 <= 1'b0;
        r_smac_hash_vld_d1 <= 1'b0;
        r_can_use_direct_path <= 1'd0;
    end else begin
        r_dmac_hash_vld_d1 <= i_dmac_hash_vld;
        r_smac_hash_vld_d1 <= i_smac_hash_vld;
        r_can_use_direct_path <= w_can_use_direct_path;
    end
end

/*======================================== �Ĵ�����ȡMAC�����???�� ========================================*/
// �Ĵ��������??����
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_reg_table_raddr <= {HASH_DATA_WIDTH{1'b0}};
    end else if (i_table_rd == 1'b1) begin
        r_reg_table_raddr <= i_table_raddr[HASH_DATA_WIDTH-1:0];
    end
end

// �Ĵ�������ʹ�ܣ��ӳ�1������RAM��ȡ??
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_reg_table_rd <= 1'b0;
    end else begin
        r_reg_table_rd <= i_table_rd;
    end
end

// ����Ĵ�����ȡ��MAC�����ݣ�ֻ�����Ч��58bit��VLAN_ID[11:0] + PORT[7:0] + MAC[47:0]??
// ��ʽ��{VLAN_ID[11:2], PORT[7:0], MAC[47:0]}
assign o_dmac_list_dout                        = { w_mac_table_rdata[VLAN_ID_WIDTH+PORT_NUM+MAC_ADDR_WIDTH-1:PORT_NUM+MAC_ADDR_WIDTH-2], 
                                                   w_mac_table_rdata[PORT_NUM+MAC_ADDR_WIDTH-1:MAC_ADDR_WIDTH], 
                                                   w_mac_table_rdata[MAC_ADDR_WIDTH-1:0]}; 

// 5������FIFO�����ݴ�����������źŷֱ�д���Ӧ��FIFO
assign w_fifo1_din = {i_vlan_id, i_rx_port};                         // VLAN_ID + RX_PORT(bitmap)
assign w_fifo2_din = i_dmac;                                         // DMAC
assign w_fifo3_din = i_smac;                                         // SMAC
assign w_fifo4_din = {i_dmac_hash_addr, i_dmac_hash_vld};            // DMAC_HASH_ADDR + DMAC_HASH_VLD
assign w_fifo5_din = {i_smac_hash_addr, i_smac_hash_vld};            // SMAC_HASH_ADDR + SMAC_HASH_VLD

// 5��FIFO��дʹ�ܣ�ͬʱд�룬ֻ�е�����FIFO������ʱ��д??
assign w_fifo1_wr_en = (w_dmac_hash_vld_posedge == 1'd1) && (w_smac_hash_vld_posedge == 1'd1) && (w_all_fifo_full == 1'd0) && (w_can_use_direct_path == 1'd0) ;
assign w_fifo2_wr_en = w_fifo1_wr_en;
assign w_fifo3_wr_en = w_fifo1_wr_en;
assign w_fifo4_wr_en = w_fifo1_wr_en;
assign w_fifo5_wr_en = w_fifo1_wr_en;

// ??5��FIFO��������н���������??
assign w_fifo_vlan_id = w_fifo1_dout[FIFO1_WIDTH-1:PORT_NUM];
assign w_fifo_rx_port = w_fifo1_dout[PORT_NUM-1:0];
assign w_fifo_dmac = w_fifo2_dout;
assign w_fifo_smac = w_fifo3_dout;
assign w_fifo_dmac_hash_addr = w_fifo4_dout[FIFO4_WIDTH-1:1];

assign w_fifo_dmac_hash_vld = w_fifo4_dout[0];
assign w_fifo_smac_hash_addr = w_fifo5_dout[FIFO5_WIDTH-1:1];

assign w_fifo_smac_hash_vld = w_fifo5_dout[0];

// 5��FIFO�Ķ�ʹ�ܣ�ͬʱ��ȡ��ֻ�е�����FIFO������ʱ�Ŷ�??
assign w_fifo1_rd_en = (r_fsm_cur_state == IDLE) && (w_all_fifo_empty == 1'd0) && (i_table_clear_req == 1'd0)  ? 1'd1 : 1'd0;
assign w_fifo2_rd_en = w_fifo1_rd_en;
assign w_fifo3_rd_en = w_fifo1_rd_en;
assign w_fifo4_rd_en = w_fifo1_rd_en;
assign w_fifo5_rd_en = w_fifo1_rd_en;

// ����FIFO����ĵ�ǰ������??
reg         [VLAN_ID_WIDTH-1:0]         r_cur_vlan_id                       ;
reg         [MAC_ADDR_WIDTH-1:0]        r_cur_dmac                          ;
reg         [HASH_DATA_WIDTH-1:0]       r_cur_dmac_hash_addr                ;       
reg         [MAC_ADDR_WIDTH-1:0]        r_cur_smac                          ;
reg         [HASH_DATA_WIDTH-1:0]       r_cur_smac_hash_addr                ;
reg         [PORT_NUM-1:0]              r_cur_rx_port                       ; // ���ն˿�bitmap

// STDģʽFIFO��ʹ���ӳټĴ���
reg                                     r_fifo_rd_en_d1                     ; // ��ʹ���ӳ�һ??

// STDģʽ��ʹ���ӳ�???��
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_fifo_rd_en_d1 <= 1'b0;
    end else begin
        r_fifo_rd_en_d1 <= w_fifo1_rd_en;
    end
end

// �ڶ�ȡFIFO��ֱ������ʱ���浱ǰ��������
// STDģʽ����rd_en����??���������ݲ���Ч������ʹ���ӳٵ�rd_en�ź� 
always @(posedge i_clk) begin
    if (i_rst) begin
        r_cur_vlan_id       <= {VLAN_ID_WIDTH{1'b0}};
        r_cur_dmac          <= {MAC_ADDR_WIDTH{1'b0}};
        r_cur_dmac_hash_addr<= {HASH_DATA_WIDTH{1'b0}};
        r_cur_smac          <= {MAC_ADDR_WIDTH{1'b0}};
        r_cur_smac_hash_addr<= {HASH_DATA_WIDTH{1'b0}};
        r_cur_rx_port       <= {PORT_NUM{1'b0}};
    end else if (r_fifo_rd_en_d1 == 1'd1) begin  // ʹ���ӳٵĶ�ʹ���ź�
        r_cur_vlan_id       <= w_fifo_vlan_id;
        r_cur_dmac          <= w_fifo_dmac;
        r_cur_dmac_hash_addr<= w_fifo_dmac_hash_addr;
        r_cur_smac          <= w_fifo_smac;
        r_cur_smac_hash_addr<= w_fifo_smac_hash_addr;
        r_cur_rx_port       <= w_fifo_rx_port;
    end else if (w_can_use_direct_path == 1'd1) begin
        r_cur_vlan_id       <= i_vlan_id;
        r_cur_dmac          <= i_dmac;
        r_cur_dmac_hash_addr<= i_dmac_hash_addr;
        r_cur_smac          <= i_smac;
        r_cur_smac_hash_addr<= i_smac_hash_addr;
        r_cur_rx_port       <= i_rx_port;
    end
end

/*---------------------------------------- 5������sync_fifoʵ��?? -------------------------------------------*/
// FIFO1: VLAN_ID + RX_PORT
sync_fifo #(
    .DEPTH                 ( INPUT_FIFO_DEPTH       ),
    .WIDTH                 ( FIFO1_WIDTH            ),
    .ALMOST_FULL_THRESHOLD ( 1                      ),
    .ALMOST_EMPTY_THRESHOLD( 1                      ),
    .FLOP_DATA_OUT         ( 0                      )  
) u_fifo1_vlan_port (
    .i_clk                 ( i_clk                  ),
    .i_rst                 ( i_rst                  ),
    .i_wr_en               ( w_fifo1_wr_en          ),
    .i_din                 ( w_fifo1_din            ),
    .o_full                ( w_fifo1_full           ),
    .i_rd_en               ( w_fifo1_rd_en          ),
    .o_dout                ( w_fifo1_dout           ),
    .o_empty               ( w_fifo1_empty          ),
    .o_almost_full         (                        ),
    .o_almost_empty        (                        ),
    .o_data_cnt            (                        )
);

// FIFO2: DMAC
sync_fifo #(
    .DEPTH                 ( INPUT_FIFO_DEPTH       ),
    .WIDTH                 ( FIFO2_WIDTH            ),
    .ALMOST_FULL_THRESHOLD ( 1                      ),
    .ALMOST_EMPTY_THRESHOLD( 1                      ),
    .FLOP_DATA_OUT         ( 0                      )  
) u_fifo2_dmac (
    .i_clk                 ( i_clk                  ),
    .i_rst                 ( i_rst                  ),
    .i_wr_en               ( w_fifo2_wr_en          ),
    .i_din                 ( w_fifo2_din            ),
    .o_full                ( w_fifo2_full           ),
    .i_rd_en               ( w_fifo2_rd_en          ),
    .o_dout                ( w_fifo2_dout           ),
    .o_empty               ( w_fifo2_empty          ),
    .o_almost_full         (                        ),
    .o_almost_empty        (                        ),
    .o_data_cnt            (                        )
);

// FIFO3: SMAC  
sync_fifo #(
    .DEPTH                 ( INPUT_FIFO_DEPTH       ),
    .WIDTH                 ( FIFO3_WIDTH            ),
    .ALMOST_FULL_THRESHOLD ( 1                      ),
    .ALMOST_EMPTY_THRESHOLD( 1                      ),
    .FLOP_DATA_OUT         ( 0                      )  
) u_fifo3_smac (
    .i_clk                 ( i_clk                  ),
    .i_rst                 ( i_rst                  ),
    .i_wr_en               ( w_fifo3_wr_en          ),
    .i_din                 ( w_fifo3_din            ),
    .o_full                ( w_fifo3_full           ),
    .i_rd_en               ( w_fifo3_rd_en          ),
    .o_dout                ( w_fifo3_dout           ),
    .o_empty               ( w_fifo3_empty          ),
    .o_almost_full         (                        ),
    .o_almost_empty        (                        ),
    .o_data_cnt            (                        )
);

// FIFO4: DMAC_HASH_ADDR + DMAC_HASH_VLD
sync_fifo #(
    .DEPTH                 ( INPUT_FIFO_DEPTH       ),
    .WIDTH                 ( FIFO4_WIDTH            ),
    .ALMOST_FULL_THRESHOLD ( 1                      ),
    .ALMOST_EMPTY_THRESHOLD( 1                      ),
    .FLOP_DATA_OUT         ( 0                      )  
) u_fifo4_dmac_hash (
    .i_clk                 ( i_clk                  ),
    .i_rst                 ( i_rst                  ),
    .i_wr_en               ( w_fifo4_wr_en          ),
    .i_din                 ( w_fifo4_din            ),
    .o_full                ( w_fifo4_full           ),
    .i_rd_en               ( w_fifo4_rd_en          ),
    .o_dout                ( w_fifo4_dout           ),
    .o_empty               ( w_fifo4_empty          ),
    .o_almost_full         (                        ),
    .o_almost_empty        (                        ),
    .o_data_cnt            (                        )
);

// FIFO5: SMAC_HASH_ADDR + SMAC_HASH_VLD
sync_fifo #(
    .DEPTH                 ( INPUT_FIFO_DEPTH       ),
    .WIDTH                 ( FIFO5_WIDTH            ),
    .ALMOST_FULL_THRESHOLD ( 1                      ),
    .ALMOST_EMPTY_THRESHOLD( 1                      ),
    .FLOP_DATA_OUT         ( 0                      )  
) u_fifo5_smac_hash (
    .i_clk                 ( i_clk                  ),
    .i_rst                 ( i_rst                  ),
    .i_wr_en               ( w_fifo5_wr_en          ),
    .i_din                 ( w_fifo5_din            ),
    .o_full                ( w_fifo5_full           ),
    .i_rd_en               ( w_fifo5_rd_en          ),
    .o_dout                ( w_fifo5_dout           ),
    .o_empty               ( w_fifo5_empty          ),
    .o_almost_full         (                        ),
    .o_almost_empty        (                        ),
    .o_data_cnt            (                        )
);

/*---------------------------------------- �����ֶν��� -------------------------------------------*/
// �����ʽ: [��Чλ[1] + �ϻ�ʱ��[AGE_TIME_WIDTH-1:0] + VLAN_ID[VLAN_ID_WIDTH-1:0] + �˿ں�[PORT_NUM-1:0] + MAC��ַ[MAC_ADDR_WIDTH-1:0]]
assign w_entry_valid    = w_mac_table_rdata[ENTRY_WIDTH-1]                                                                    ;
assign w_entry_age_time = w_mac_table_rdata[ENTRY_WIDTH-2:ENTRY_WIDTH-1-AGE_TIME_WIDTH]                                       ;  
assign w_entry_vlan_id  = w_mac_table_rdata[ENTRY_WIDTH-1-AGE_TIME_WIDTH-1:ENTRY_WIDTH-1-AGE_TIME_WIDTH-VLAN_ID_WIDTH]        ;
assign w_entry_port     = w_mac_table_rdata[PORT_NUM+MAC_ADDR_WIDTH-1:MAC_ADDR_WIDTH]                                         ;
assign w_entry_mac      = w_mac_table_rdata[MAC_ADDR_WIDTH-1:0]                                                               ;

/*---------------------------------------- bitmap��Ч�Լ�?? ----------------------------------------------*/
// ??��r_cur_rx_port�Ƿ�Ϊ��Ч��one-hot����(ֻ��??��bit??1)��ȫ0
wire                                    w_rx_port_valid                     ; // ���ն˿�bitmap��Ч��־
wire  [AGE_TIME_WIDTH-1:0]              w_age_time_diff                     ;
assign w_rx_port_valid = (r_cur_rx_port != {PORT_NUM{1'b0}}) && ((r_cur_rx_port & (r_cur_rx_port - {{(PORT_NUM-1){1'b0}}, 1'b1})) == {PORT_NUM{1'b0}}) ? 1'd1 : 1'd0;

/*---------------------------------------- ƥ���߼� ----------------------------------------------*/
assign w_dmac_match     = (w_entry_valid == 1'd1 && (w_entry_mac == r_cur_dmac) && (w_entry_vlan_id == r_cur_vlan_id)) ? 1'd1 : 1'd0      ;
assign w_smac_match     = (w_entry_valid == 1'd1 && (w_entry_mac == r_cur_smac) && (w_entry_vlan_id == r_cur_vlan_id)) ? 1'd1 : 1'd0      ;
assign w_smac_port_match= (w_smac_match  == 1'd1 && w_rx_port_valid == 1'd1 && (w_entry_port == r_cur_rx_port)) ? 1'd1 : 1'd0 ;

// �ϻ�??��???��??  ��ǰʱ�����ȥ����ʱ����Ĳ�ֵ���ڵ���???����???ʱ��Ϊ����
assign w_entry_expired  = w_entry_valid == 1'd1 && (r_entry_expired_flag == 1'd1) ? 1'd1 : 1'd0 ;
assign w_age_time_diff = r_global_timestamp - w_entry_age_time;
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_entry_expired_flag <= 1'b0;
    end else begin
        r_entry_expired_flag <= (w_age_time_diff >= i_age_time_threshold) && w_entry_valid == 1'd1 ? 1'd1 : 1'd0;
    end
end
/*---------------------------------------- ����??��???�� -------------------------------------------*/
assign w_table_full     = (r_table_entry_cnt >= i_table_full_threshold) ? 1'd1 : 1'd0                   ;

always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_table_full <= 1'b0;
    end else begin
        r_table_full <= w_table_full;
    end
end

always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_dmac_list_full_er_stat <= 1'b0;
    end else if (i_table_clear_req) begin
        r_dmac_list_full_er_stat <= 1'b0;
    end else begin
        r_dmac_list_full_er_stat <= w_table_full == 1'b1 && r_table_full == 1'b0 ? 1'b1 : 1'b0;
    end
end

always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_dmac_list_full_er_cnt <= 16'd0;
    end else if (i_table_clear_req) begin
        r_dmac_list_full_er_cnt <= 16'd0;
    end else begin
        r_dmac_list_full_er_cnt <= w_table_full == 1'b1 && r_table_full == 1'b0 ? r_dmac_list_full_er_cnt + 1'd1 : r_dmac_list_full_er_cnt;
    end
end

/*---------------------------------------- �ϻ�ɨ�败���߼� -------------------------------------------*/
// 32bit�ֳ�4�αȽϣ�ÿ��8bit
wire w_age_scan_flag0 ;
wire w_age_scan_flag1 ;
wire w_age_scan_flag2 ;
wire w_age_scan_flag3 ;

assign w_age_scan_flag0 = (r_age_scan_timer[7:0]   >= i_age_scan_interval[7:0]);
assign w_age_scan_flag1 = (r_age_scan_timer[15:8]  >= i_age_scan_interval[15:8]);
assign w_age_scan_flag2 = (r_age_scan_timer[23:16] >= i_age_scan_interval[23:16]);
assign w_age_scan_flag3 = (r_age_scan_timer[31:24] >= i_age_scan_interval[31:24]);

assign w_age_scan_trigger = (w_age_scan_flag0 == 1'd1 && w_age_scan_flag1 == 1'd1 && w_age_scan_flag2 == 1'd1 && w_age_scan_flag3 == 1'd1) && (r_table_entry_cnt > 15'd0) ? 1'd1 : 1'd0;

/*---------------------------------------- �����??? -------------------------------------------*/
assign o_dmac_lookup_vld    = r_dmac_lookup_vld                                                           ;
assign o_dmac_tx_port       = r_dmac_tx_port                                                              ;
assign o_dmac_lookup_hit    = r_dmac_lookup_hit                                                           ;
assign o_lookup_clash       = r_lookup_clash                                                              ;
assign o_table_full         = w_table_full                                                                ;
//assign o_reg_bus_rdata      = r_reg_bus_rdata                                                             ;
//assign o_reg_bus_rdata_vld  = r_reg_bus_rdata_vld                                                         ;


/*======================================== ״???��  ========================================*/
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_fsm_cur_state <= IDLE;
    end else begin
        r_fsm_cur_state <= r_fsm_nxt_state;
    end
end

always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_state_cnt <= 16'd0;
    end else if (r_fsm_cur_state != r_fsm_nxt_state) begin
        r_state_cnt <= 16'd0;
    end else begin
        r_state_cnt <= r_state_cnt + 1'b1;  
    end
end

always @(*) begin
    r_fsm_nxt_state = r_fsm_cur_state;   
    case (r_fsm_cur_state)
        IDLE: 
            r_fsm_nxt_state = (i_table_clear_req == 1'd1) ? AGE_SCAN :       // ������ȼ���??
                              // ??��FIFO�Ƿ������ݿɴ������ֱ�����ݿ���
                              (r_can_use_direct_path == 1'd1) ? DMAC_LOOKUP :  // ֱ��·�������ȴ�״???
                              (w_all_fifo_empty == 1'd0) ? FIFO_READ_WAIT :    // STDģʽ??Ҫ�ȴ�����׼??
                              (r_age_scan_en == 1'd1) ? AGE_SCAN :             // �ϻ�ɨ��
                              IDLE;
        FIFO_READ_WAIT:   // STDģʽFIFO��ȡ�ȴ�״???
            r_fsm_nxt_state = DMAC_LOOKUP;                                    // �ȴ�??�����ں�����׼���ã�������
        DMAC_LOOKUP:   
            r_fsm_nxt_state = (r_state_cnt == 16'd1 &&  w_dmac_match == 1'd1) ? DMAC_REFRESH :  
                              (r_state_cnt == 16'd1 &&  w_dmac_match == 1'd0) ? SMAC_LEARN_CHECK : DMAC_LOOKUP;// ƥ����ˢ��???��ʱ�� ��Ȼ��ѧϰSMAC                                          
        DMAC_REFRESH: 
            r_fsm_nxt_state = SMAC_LEARN_CHECK;                     // ˢ����ɣ�����SMACѧϰ        
        SMAC_LEARN_CHECK: 
            r_fsm_nxt_state = ((w_smac_match == 1'd1) || ((w_entry_valid == 1'd0) && (w_table_full == 1'd0))) ? SMAC_LEARN_UPDATE :  // SMAC+VLANƥ���ձ����ѧ??
                              IDLE;                                  // ��ϣ��ͻ��MAC+VLAN��ƥ�䣩������������ؿ�??        
        SMAC_LEARN_UPDATE: 
            r_fsm_nxt_state = (r_state_cnt == 16'd1) ? IDLE : SMAC_LEARN_UPDATE;   // �ȴ�1��ʱ��������RAM�����ȶ��󷵻�IDLE        
        AGE_SCAN: 
            r_fsm_nxt_state = (r_mac_table_addr == {HASH_DATA_WIDTH{1'b1}}) ? IDLE :    // ɨ����ɣ����������ɣ�
                              ((w_new_packet_arrival == 1'd1) && ((i_table_clear_req == 1'd0) || (r_clear_burst_cnt >= CLEAR_BURST_LIMIT))) ? IDLE : // �б��ĵȴ���(�����ģ?? ?? �Ѵﵽͻ����??)ʱ�����ȴ�����
                              ((w_entry_valid == 1'd1) && (w_entry_expired == 1'd1) && (i_table_clear_req == 1'd0) && (r_state_cnt >= 16'd1)) ? AGE_UPDATE :    // ??Ҫ???�����£������ģʽ����ȷ�������ȶ�
                              AGE_SCAN;                                              // ����ɨ����һ����??        
        AGE_UPDATE: 
            r_fsm_nxt_state = (r_mac_table_addr == {HASH_DATA_WIDTH{1'b1}}) ? IDLE :  // ɨ�����
                              ((w_all_fifo_empty == 1'd0) && ((i_table_clear_req == 1'd0) || (r_clear_burst_cnt >= CLEAR_BURST_LIMIT))) ? IDLE : // �б��ĵȴ���(�����ģ?? ?? �Ѵﵽͻ����??)ʱ�����ȴ�����
                              AGE_SCAN;                                                // �ϻ�������ɣ�����ɨ??        
        default: 
            r_fsm_nxt_state = IDLE;
    endcase
end

/*========================================  �������ݹ��� ========================================*/
/*
// FIFO���뻺�����֧����������???���Ḳ�����ڴ��������
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_reg_bus_we          <= 1'b0;
        r_reg_bus_addr        <= {REG_ADDR_BUS_WIDTH{1'b0}};
        r_reg_bus_data        <= {REG_DATA_BUS_WIDTH{1'b0}};
        r_reg_bus_data_vld    <= 1'b0;
        r_reg_bus_re          <= 1'b0;
        r_reg_bus_raddr       <= {REG_ADDR_BUS_WIDTH{1'b0}};
    end else begin
        r_reg_bus_we       <= i_reg_bus_we;
        r_reg_bus_addr     <= i_reg_bus_addr;
        r_reg_bus_data     <= i_reg_bus_data;
        r_reg_bus_data_vld <= i_reg_bus_data_vld;
        r_reg_bus_re       <= i_reg_bus_re;
        r_reg_bus_raddr    <= i_reg_bus_raddr;
    end
end
*/
/*======================================== ���üĴ�����?? ========================================*/
/*
// �ϻ�ʱ����???���üĴ���
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_age_time_threshold <= 10'd300;
    end else if(SIM_MODE == 1) begin
        r_age_time_threshold <= 10'd8;
    end else if ((r_reg_bus_we == 1'd1) && (r_reg_bus_data_vld == 1'd1) && (r_reg_bus_addr == REG_AGE_TIME_THRESHOLD)) begin
        r_age_time_threshold <= r_reg_bus_data[AGE_TIME_WIDTH-1:0];
    end
end

// ���������Ĵ���
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_table_clear_req <= 1'b0;
    end else if ((r_reg_bus_we == 1'd1) && (r_reg_bus_data_vld == 1'd1) && (r_reg_bus_addr == REG_TABLE_CLEAR)) begin
        r_table_clear_req <= r_reg_bus_data[0];
    end else if ((r_table_clear_req == 1'd1) && (r_mac_table_addr == {HASH_DATA_WIDTH{1'b1}}) && (r_fsm_cur_state == AGE_SCAN)) begin
        r_table_clear_req <= 1'b0;
    end
end

// ������???���üĴ���
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_table_full_threshold <= TABLE_FULL_THRESHOLD;
    end else if ((r_reg_bus_we == 1'd1) && (r_reg_bus_data_vld == 1'd1) && (r_reg_bus_addr == REG_TABLE_FULL_THRESHOLD)) begin
        r_table_full_threshold <= r_reg_bus_data[14:0];
    end
end

// �ϻ�ɨ�������üĴ�??
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_age_scan_interval <= AGE_SCAN_INTERVAL;
    end else if ((r_reg_bus_we == 1'd1) && (r_reg_bus_data_vld == 1'd1) && (r_reg_bus_addr == REG_AGE_SCAN_INTERVAL)) begin
        r_age_scan_interval <= {{16{1'b0}}, r_reg_bus_data};
    end
end
*/
/*======================================== ͳ�Ƽ�������?? ========================================*/
// MACѧϰ�ɹ�ͳ�Ƽ���??  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_learn_success_cnt <= 32'd0;
    end else if (i_table_clear_req == 1'd1) begin
        r_learn_success_cnt <= 32'd0;
    end else if ((r_fsm_cur_state == SMAC_LEARN_UPDATE) && (r_state_cnt == 16'd1)) begin
        if ((w_smac_match == 1'd1) || ((w_entry_valid == 1'd0) && w_rx_port_valid == 1'd1 && (w_table_full == 1'd0))) begin
            r_learn_success_cnt <= r_learn_success_cnt + 1'b1;
        end
    end
end

// MACѧϰʧ��ͳ�Ƽ���??  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_learn_fail_cnt <= 32'd0;
    end else if (i_table_clear_req == 1'd1) begin
        r_learn_fail_cnt <= 32'd0;
    end else if ((r_fsm_cur_state == SMAC_LEARN_UPDATE) && (r_state_cnt == 16'd1)) begin
        if (((w_entry_valid == 1'd1) && (w_smac_match == 1'd0)) || ((w_entry_valid == 1'd0) && (w_table_full == 1'd1)) || (w_rx_port_valid == 1'd0)) begin
            r_learn_fail_cnt <= r_learn_fail_cnt + 1'b1;
        end
    end else if (r_fsm_cur_state == SMAC_LEARN_CHECK) begin
        if ((w_entry_valid == 1'd0) && (w_table_full == 1'd1)) begin
            r_learn_fail_cnt <= r_learn_fail_cnt + 1'b1;
        end
    end
end

// ��ϣ��ͻͳ�Ƽ���??  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_collision_cnt <= 32'd0;
    end else if (i_table_clear_req) begin
        r_collision_cnt <= 32'd0;
    end else if (r_fsm_cur_state == DMAC_LOOKUP && r_state_cnt == 16'd1 && w_entry_valid == 1'd1 && w_dmac_match == 1'd0) begin
        r_collision_cnt <= r_collision_cnt + 1'b1;
    end else if (r_fsm_cur_state == SMAC_LEARN_UPDATE && r_state_cnt == 16'd1 && w_entry_valid == 1'd1 && w_smac_match == 1'd0) begin
        r_collision_cnt <= r_collision_cnt + 1'b1;
    end
end

// �˿��ƶ�ͳ�Ƽ���??  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_port_move_cnt <= 32'd0;
    end else if (i_table_clear_req) begin
        r_port_move_cnt <= 32'd0;
    end else if (r_fsm_cur_state == SMAC_LEARN_UPDATE && r_state_cnt == 16'd1) begin
        if (w_smac_match == 1'd1 && w_rx_port_valid == 1'd1 && (w_entry_port != r_cur_rx_port)) begin
            r_port_move_cnt <= r_port_move_cnt + 1'b1;
        end
    end
end

/*======================================== �����������?? ========================================*/
// �������?? - ������ЧMAC������������ֹ���������
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_table_entry_cnt <= 15'd0;
    end else if (i_table_clear_req) begin
        r_table_entry_cnt <= 15'd0;
    end else if (r_entry_add == 1'd1 && r_entry_del == 1'd0) begin
        if (r_table_entry_cnt < 15'h7FFF) begin  
            r_table_entry_cnt <= r_table_entry_cnt + 1'b1;  
        end
    end else if (r_entry_add == 1'd0 && r_entry_del == 1'd1) begin
        if (r_table_entry_cnt > 15'd0) begin  
            r_table_entry_cnt <= r_table_entry_cnt - 1'b1; 
        end
    end
end

/*======================================== �Ĵ����������߼� ========================================*/
// �Ĵ����������߼�
/*
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_reg_bus_rdata <= {REG_DATA_BUS_WIDTH{1'b0}};
    end else if (r_reg_bus_re) begin
        case (r_reg_bus_raddr)
            REG_AGE_TIME_THRESHOLD: begin
                // ��???Ӧλ��:ֱ�ӽ�ȡ����??,��ֹREG_DATA_BUS_WIDTH<AGE_TIME_WIDTHʱ��??
                r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_age_time_threshold[AGE_TIME_WIDTH-1:0];
            end
            REG_TABLE_CLEAR: begin
                r_reg_bus_rdata <= {{(REG_DATA_BUS_WIDTH-1){1'b0}}, r_table_clear_req};
            end
            REG_TABLE_FULL_THRESHOLD: begin
                // ��???Ӧλ��:ֱ�ӽ�ȡ��λ,��ֹREG_DATA_BUS_WIDTH<15ʱ��??
                r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_table_full_threshold[14:0];
            end
            REG_AGE_SCAN_INTERVAL: begin 
                r_reg_bus_rdata <= r_age_scan_interval[REG_DATA_BUS_WIDTH-1:0]; 
            end
            REG_TABLE_ENTRY_cnt: begin 
                // ��???Ӧλ��:ֱ�ӽ�ȡ��λ,��ֹREG_DATA_BUS_WIDTH<15ʱ��??
                r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_table_entry_cnt[14:0]; 
            end
            REG_LEARN_STATISTICS: begin
                r_reg_bus_rdata <= {r_learn_success_cnt[15:0]};
            end
            REG_COLLISION_STATISTICS: begin
                r_reg_bus_rdata <= r_collision_cnt[REG_DATA_BUS_WIDTH-1:0];
            end
            REG_PORT_MOVE_STATISTICS: begin
                r_reg_bus_rdata <= r_port_move_cnt[REG_DATA_BUS_WIDTH-1:0];
            end
            default: begin
                r_reg_bus_rdata <= {REG_DATA_BUS_WIDTH{1'b0}};
            end
        endcase
    end else begin
        r_reg_bus_rdata <= {REG_DATA_BUS_WIDTH{1'b0}};
    end
end
// �Ĵ�����������Ч��־
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_reg_bus_rdata_vld <= 1'b0;
    end else begin
        r_reg_bus_rdata_vld <= r_reg_bus_re;
    end
end
*/
/*======================================== ʱ�����?? ========================================*/
// ΢�����??  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_us_cnt <= 16'd0;
    end else if (r_us_cnt >= US_CNT_MAX - 1) begin
        r_us_cnt <= 16'd0;
    end else begin
        r_us_cnt <= r_us_cnt + 1'b1;
    end
end

// ΢�������ź�����  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_us_pulse <= 1'b0;
    end else begin
        r_us_pulse <= (r_us_cnt == US_CNT_MAX - 1);
    end
end
// �������??  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_ms_cnt <= 10'd0;
    end else if (r_us_pulse) begin
        if (r_ms_cnt >= MS_CNT_MAX - 1) begin
            r_ms_cnt <= 10'd0;
        end else begin
            r_ms_cnt <= r_ms_cnt + 1'b1;
        end
    end
end

// ���������ź�����  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_ms_pulse <= 1'b0;
    end else begin
        r_ms_pulse <= r_us_pulse == 1'd1 && (r_ms_cnt == MS_CNT_MAX - 1) ? 1'd1 : 1'd0;
    end
end

// �����ܼ����� 
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_s_cnt <= 32'd0;
    end else if (r_ms_pulse) begin
        if (r_s_cnt >= S_CNT_MAX - 1) begin
            r_s_cnt <= 32'd0;
        end else begin
            r_s_cnt <= r_s_cnt + 1'b1;
        end
    end
end

// 1�������ź���??  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_age_timer_pulse <= 1'b0;
    end else begin
        r_age_timer_pulse <= r_ms_pulse == 1'd1 && (r_s_cnt == S_CNT_MAX - 1) ? 1'd1 : 1'd0;
    end
end

// ȫ��ʱ���������  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_global_timestamp <= {AGE_TIME_WIDTH{1'b0}};
    end else if (r_age_timer_pulse) begin
        r_global_timestamp <= r_global_timestamp + 1'b1;
    end
end

// �ϻ�ɨ��������??
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_age_scan_timer <= 32'd0;
    end else if (w_age_scan_trigger) begin
        r_age_scan_timer <= 32'd0;
    end else if (r_age_timer_pulse == 1'd1 && r_table_entry_cnt > 15'd0) begin
        r_age_scan_timer <= r_age_scan_timer + 1'b1;
    end
end

/*======================================== ���ͻ�������߼� ========================================*/
// ���ͻ������?? 
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_clear_burst_cnt <= 8'd0;
    end else if (r_fsm_cur_state != AGE_SCAN || i_table_clear_req == 1'd0) begin
        r_clear_burst_cnt <= 8'd0;
    end else if (r_fsm_cur_state == AGE_SCAN && i_table_clear_req == 1'd1) begin
        if (r_clear_burst_cnt < CLEAR_BURST_LIMIT) begin
            r_clear_burst_cnt <= r_clear_burst_cnt + 1'b1;
        end
    end
end

/*======================================== �ϻ�ɨ���ַ���� ========================================*/
// �ϻ�ɨ��ϵ��ַ����
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_age_scan_breakpoint <= {HASH_DATA_WIDTH{1'b0}};
    end else if (r_fsm_cur_state == AGE_SCAN && r_fsm_nxt_state == IDLE && r_mac_table_addr != {HASH_DATA_WIDTH{1'b1}}) begin
        r_age_scan_breakpoint <= r_mac_table_addr;  // �����ʱ���浱ǰ��ַ
    end else if (r_mac_table_addr == {HASH_DATA_WIDTH{1'b1}}) begin
        r_age_scan_breakpoint <= {HASH_DATA_WIDTH{1'b0}};  // ɨ�����ʱ���ö�??
    end
end

// �ϻ�ɨ��ʹ���ź� 
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_age_scan_en <= 1'b0;
    end else if (r_mac_table_addr == {HASH_DATA_WIDTH{1'b1}}) begin
        r_age_scan_en <= 1'b0;
    end else if (w_age_scan_trigger) begin
        r_age_scan_en <= 1'b1;
    end
end

/*======================================== MAC��洢�����ʿ��� ========================================*/
// MAC���??����  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_mac_table_addr <= {HASH_DATA_WIDTH{1'b0}};
    end else begin
        case (r_fsm_cur_state)
            IDLE: begin
                if (r_can_use_direct_path == 1'd1||w_can_use_direct_path == 1'd1) begin
                    r_mac_table_addr <= i_dmac_hash_addr;  // ֱ��·����������ʹ��
                end else if (w_all_fifo_empty == 1'd0) begin
                    // STDģʽ����������ʹ��FIFO�������Ҫ�ȶ�ȡ������FIFO_READ_WAIT״???��??
                    r_mac_table_addr <= {HASH_DATA_WIDTH{1'b0}};  // ����??
                end else begin
                    r_mac_table_addr <= {HASH_DATA_WIDTH{1'b0}};
                end
            end
            FIFO_READ_WAIT: begin  // �ڴ�״???���ô����������л�ȡ�ĵ�ַ
                r_mac_table_addr <= r_cur_dmac_hash_addr;  // ʹ�������������
            end
            DMAC_LOOKUP: begin 
                r_mac_table_addr <= r_state_cnt == 16'd1 &&  w_dmac_match == 1'd0 ? r_cur_smac_hash_addr : r_cur_dmac_hash_addr;  // ʹ�������������
            end
            DMAC_REFRESH: begin
                r_mac_table_addr <= r_cur_smac_hash_addr;
            end
            SMAC_LEARN_CHECK, SMAC_LEARN_UPDATE: begin
                r_mac_table_addr <= r_cur_smac_hash_addr;
            end
            AGE_SCAN, AGE_UPDATE: begin
                if (r_fsm_cur_state == IDLE && (r_fsm_nxt_state == AGE_SCAN)) begin
                    r_mac_table_addr <= r_age_scan_breakpoint;  // �Ӷϵ�ָ���??0????
                end else if (r_fsm_cur_state == AGE_SCAN) begin
                    if (i_table_clear_req == 1'd1) begin
                        if (r_mac_table_addr != {HASH_DATA_WIDTH{1'b1}}) begin
                            r_mac_table_addr <= r_mac_table_addr + 1'b1;
                        end
                    end else begin
                        if (r_fsm_nxt_state == AGE_UPDATE) begin
                            r_mac_table_addr <= r_mac_table_addr;
                        end else if ((r_mac_table_addr != {HASH_DATA_WIDTH{1'b1}}) && (r_agescan_cnt == 1'd1)) begin
                            r_mac_table_addr <= r_mac_table_addr + 1'b1;
                        end
                    end
                end else if (r_fsm_cur_state == AGE_UPDATE) begin
                    if (r_fsm_nxt_state == AGE_SCAN) begin
                        if (r_mac_table_addr != {HASH_DATA_WIDTH{1'b1}}) begin
                            r_mac_table_addr <= r_mac_table_addr + 1'b1;
                        end
                    end else begin
                        r_mac_table_addr <= r_mac_table_addr;
                    end
                end
            end
            default: begin
                r_mac_table_addr <= {HASH_DATA_WIDTH{1'b0}};
            end
        endcase
    end
end

// ��AGE_SCNAʱ����ַ״???������??
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_agescan_cnt <= 1'd0;
    end else if (r_mac_table_re == 1'd1 && r_fsm_cur_state == AGE_SCAN) begin
        r_agescan_cnt <= r_agescan_cnt == 1'd0 ? 1'd1 : 1'd0;
    end else begin
        r_agescan_cnt <= 1'd0;
    end
end

// MAC���ʹ�ܿ���  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_mac_table_re <= 1'b0;
    end else begin
        case (r_fsm_cur_state)
            IDLE: begin
                r_mac_table_re <= ((r_can_use_direct_path == 1'd1||w_can_use_direct_path == 1'd1) || (w_all_fifo_empty == 1'd0)) && (i_table_clear_req == 1'd0) ? 1'd1 : 1'd0;
            end
            FIFO_READ_WAIT: begin  // FIFO��ȡ�ȴ�״???������RAM��ȡ
                r_mac_table_re <= 1'b1;
            end
            DMAC_LOOKUP, SMAC_LEARN_CHECK: begin
                r_mac_table_re <= 1'b1;
            end
            DMAC_REFRESH: begin
                r_mac_table_re <= 1'b0;
            end
            SMAC_LEARN_UPDATE: begin
                r_mac_table_re <= 1'b0;
            end
            AGE_SCAN: begin
                if ((i_table_clear_req == 1'd1) && (r_fsm_nxt_state == AGE_UPDATE)) begin
                    r_mac_table_re <= 1'b0;
                end else if(((r_state_cnt == 1'd0) || !((w_entry_valid == 1'd1) && (w_entry_expired == 1'd1)))  )begin
                    r_mac_table_re <= 1'b1;
                end else begin
                    r_mac_table_re <= 1'b0;
                end
            end
            AGE_UPDATE: begin
                r_mac_table_re <= 1'b1;
            end
            default: begin
                r_mac_table_re <= 1'b0;
            end
        endcase
    end
end

// MAC��дʹ�ܿ���  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_mac_table_we <= 1'b0;
    end else begin
        case (r_fsm_cur_state)
            DMAC_REFRESH: begin
                r_mac_table_we <= 1'b1;
            end
            SMAC_LEARN_UPDATE: begin
                if (r_state_cnt == 16'd1) begin
                    r_mac_table_we <= (w_smac_match || (w_entry_valid == 1'd0 && w_rx_port_valid == 1'd1 && w_table_full == 1'd0));
                end else begin
                    r_mac_table_we <= 1'b0;  
                end
            end
            AGE_SCAN: begin
                if (i_table_clear_req) begin
                    r_mac_table_we <= 1'b1;
                end else begin
                    r_mac_table_we <= r_fsm_nxt_state == AGE_UPDATE ? 1'b1 : 1'b0;
                end
            end
            AGE_UPDATE: begin
                r_mac_table_we <= 1'b0;
            end
            default: begin
                r_mac_table_we <= 1'b0;
            end
        endcase
    end
end

// MAC��д���ݿ��� - ʹ�õ�ǰ����Ļ�����??
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_mac_table_wdata <= {ENTRY_WIDTH{1'b0}};
    end else begin
        case (r_fsm_cur_state)
            DMAC_REFRESH: begin
                r_mac_table_wdata <= {w_entry_valid, r_global_timestamp, w_entry_vlan_id, 
                                    w_entry_port, w_entry_mac};
            end
            SMAC_LEARN_UPDATE: begin
                if (r_state_cnt == 16'd1) begin
                    if (w_smac_match) begin
                        if (w_smac_port_match) begin
                            r_mac_table_wdata <= {1'b1, r_global_timestamp, w_entry_vlan_id, 
                                                w_entry_port, w_entry_mac};
                        end else begin
                            r_mac_table_wdata <= {1'b1, 
                                                r_global_timestamp[AGE_TIME_WIDTH-1:0], 
                                                r_cur_vlan_id[VLAN_ID_WIDTH-1:0], 
                                                r_cur_rx_port[PORT_NUM-1:0], 
                                                r_cur_smac[MAC_ADDR_WIDTH-1:0]};
                        end
                    end else if (w_entry_valid == 1'd0 && w_rx_port_valid == 1'd1 && w_table_full == 1'd0) begin
                        r_mac_table_wdata <= {1'b1, 
                                            r_global_timestamp[AGE_TIME_WIDTH-1:0], 
                                            r_cur_vlan_id[VLAN_ID_WIDTH-1:0], 
                                            r_cur_rx_port[PORT_NUM-1:0], 
                                            r_cur_smac[MAC_ADDR_WIDTH-1:0]};
                    end else begin  
                        r_mac_table_wdata <= w_mac_table_rdata;
                    end
                end else begin
                    r_mac_table_wdata <= r_mac_table_wdata;
                end
            end
            AGE_UPDATE: begin
                r_mac_table_wdata <= {ENTRY_WIDTH{1'b0}};
            end
            AGE_SCAN: begin
                if (i_table_clear_req) begin
                    r_mac_table_wdata <= {ENTRY_WIDTH{1'b0}};
                end else if (w_entry_valid == 1'd1 && w_entry_expired == 1'd1) begin
                    r_mac_table_wdata <= {ENTRY_WIDTH{1'b0}};
                end else begin
                    r_mac_table_wdata <= w_mac_table_rdata; 
                end
            end
            default: begin
                r_mac_table_wdata <= {ENTRY_WIDTH{1'b0}};
            end
        endcase
    end
end

/*======================================== ������������߼� ========================================*/
// ������ӱ�־����  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_entry_add <= 1'b0;
    end else if (r_fsm_cur_state == SMAC_LEARN_UPDATE && r_state_cnt == 16'd1 && 
                 w_entry_valid == 1'd0 && w_rx_port_valid == 1'd1 && w_table_full == 1'd0) begin
        r_entry_add <= 1'b1;
    end else begin
        r_entry_add <= 1'b0;
    end
end

// ����ɾ����־����  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_entry_del <= 1'b0;
    end else if (r_fsm_cur_state == AGE_UPDATE && w_entry_valid == 1'd1 && w_entry_expired == 1'd1) begin
        r_entry_del <= 1'b1;
    end else if (r_fsm_cur_state == AGE_SCAN && i_table_clear_req == 1'd1 && w_entry_valid == 1'd1) begin
        r_entry_del <= 1'b1;
    end else begin
        r_entry_del <= 1'b0;
    end
end

/*======================================== ��������߼� ========================================*/
// DMAC�������Ч��־  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_dmac_lookup_vld <= 1'b0;
    end else if (r_fsm_cur_state == DMAC_LOOKUP && r_state_cnt == 16'd1) begin
        r_dmac_lookup_vld <= 1'b1;
    end else begin
        r_dmac_lookup_vld <= 1'b0;
    end
end

// DMAC������б�־  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_dmac_lookup_hit <= 1'b0;
    end else if (r_fsm_cur_state == DMAC_LOOKUP && r_state_cnt == 16'd1) begin
        r_dmac_lookup_hit <= w_dmac_match;
    end else begin
        r_dmac_lookup_hit <= 1'b0;
    end
end

// DMACת���˿�  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_dmac_tx_port <= {PORT_NUM{1'b0}};
    end else if (r_fsm_cur_state == DMAC_LOOKUP && r_state_cnt == 16'd1) begin
        if (w_dmac_match) begin
            r_dmac_tx_port <= w_entry_port;
        end else begin
            r_dmac_tx_port <= {PORT_NUM{1'b0}};  // δ�鵽ʱֱ�����0
        end
    end else begin
        r_dmac_tx_port <= {PORT_NUM{1'b0}};
    end
end

// ����ͻ??��???��  
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_lookup_clash <= 1'b0;
    end else if (r_fsm_cur_state == DMAC_LOOKUP && r_state_cnt == 16'd1) begin
        r_lookup_clash <= w_entry_valid == 1'd1 && w_dmac_match == 1'd0;
    end else begin
        r_lookup_clash <= 1'b0;
    end
end

/*======================================== MAC���?? ========================================*/

ram_simple2port #(
    .RAM_WIDTH      ( ENTRY_WIDTH               ),
    .RAM_DEPTH      ( MAC_TABLE_DEPTH           ),
    .RAM_PERFORMANCE( "LOW_LATENCY"             ), 
    .INIT_FILE      (  0                        )  
) u_mac_table_ram (
    .addra          ( r_mac_table_addr                      ),
    .addrb          ( r_mac_table_addr                      ),
    .dina           ( r_mac_table_wdata                     ), 
    .clka           ( i_clk                                 ), 
    .clkb           ( i_clk                                 ), 
    .wea            ( r_mac_table_we                        ), // ѧϰ
    .enb            ( r_mac_table_re                        ), // ���
    .rstb           ( i_rst                                 ), 
    .regceb         ( 1'b0                                  ),
    .doutb          ( w_mac_table_rdata                     )  
);

endmodule