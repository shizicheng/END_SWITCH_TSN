module rx_mac_hash_calc#(  
    parameter           CWIDTH              =           15
)(
    input               wire                                    i_clk                   ,   // 250MHz
    input               wire                                    i_rst                   ,
    /*---------------------------------------- �Ĵ������ýӿ� -------------------------------------------*/
    input               wire   [15:0]                           i_hash_poly_regs        ,
    input               wire   [15:0]                           i_hash_init_val_regs    ,
    input               wire                                    i_hash_regs_vld         ,
    /*--------------------------------- ��Ϣ��ȡģ������� MAC ��Ϣ -------------------------------------*/
    input               wire   [11:0]                           i_vlan_id               , // ���뱨�ĵ�VLAN ID
    input               wire   [47:0]                           i_dmac_data             , // Ŀ�� MAC ��ַ(48bit)
    input               wire                                    i_dmac_data_vld         , // DMAC������Ч
    input               wire   [47:0]                           i_smac_data             , // Դ MAC ��ַ(48bit)
    input               wire                                    i_smac_data_vld         , // SMAC������Ч
    /*--------------------------------- ��� hash �ļ����� -------------------------------------*/     
    output              wire   [11:0]                           o_vlan_id               ,
    output              wire   [CWIDTH - 1 : 0]                 o_dmac_hash_key         ,
    output              wire   [47 : 0]                         o_dmac                  ,
    output              wire                                    o_dmac_hash_vld         , 
    output              wire   [CWIDTH - 1 : 0]                 o_smac_hash_key         ,
    output              wire   [47 : 0]                         o_smac                  ,
    output              wire                                    o_smac_hash_vld               
);

// �����źŴ���
reg     [47:0]                              ri_dmac_data                        ; // DMAC ���ݴ���(48bit)
reg                                         ri_dmac_data_vld                    ; // DMAC ������Ч����
reg     [47:0]                              ri_smac_data                        ; // SMAC ���ݴ���(48bit)
reg                                         ri_smac_data_vld                    ; // SMAC ������Ч����
reg     [11:0]                              ri_vlan_id                          ; // VLAN ID����

// �ڲ��������
reg                                         r_dmac_hash_en                      ; // DMAC HASH ʹ��
reg                                         r_smac_hash_en                      ; // SMAC HASH ʹ��
reg                                         r_dmac_hash_vld                     ; // DMAC HASH ��Ч
reg                                         r_smac_hash_vld                     ; // SMAC HASH ��Ч

// ����Ĵ���
reg     [11:0]                              ro_vlan_id                          ; // VLAN ID ���
reg     [CWIDTH-1:0]                        ro_dmac_hash_key                    ; // DMAC HASH KEY ���
reg     [47:0]                              ro_dmac                             ; // DMAC ���
// reg                                         ro_dmac_vld                         ; // DMAC ��Ч���
reg     [CWIDTH-1:0]                        ro_smac_hash_key                    ; // SMAC HASH KEY ���
reg     [47:0]                              ro_smac                             ; // SMAC ���
// reg                                         ro_smac_vld                         ; // SMAC ��Ч���
reg                                         r_hash_cacl_rst                     ;

// HASH �������
wire    [CWIDTH-1:0]                        w_dmac_crc_out                      ; // DMAC CRC ���
wire    [CWIDTH-1:0]                        w_smac_crc_out                      ; // SMAC CRC ���

//---------- ����źŸ�ֵ ----------
assign  o_vlan_id                           =       ro_vlan_id                  ;
assign  o_dmac_hash_key                     =       ro_dmac_hash_key            ;
assign  o_dmac                              =       ro_dmac                     ;
assign  o_dmac_hash_vld                     =       r_dmac_hash_vld             ;
assign  o_smac_hash_key                     =       ro_smac_hash_key            ;
assign  o_smac                              =       ro_smac                     ;
assign  o_smac_hash_vld                     =       r_smac_hash_vld             ;
 
// �����źŴ���
always @(posedge i_clk) begin
    if (i_rst) begin
        ri_dmac_data     <= 48'd0;
        ri_dmac_data_vld <= 1'b0;
        ri_smac_data     <= 48'd0;
        ri_smac_data_vld <= 1'b0;
        ri_vlan_id       <= 12'd0;
    end else begin
        ri_dmac_data     <= i_dmac_data_vld ? i_dmac_data : ri_dmac_data;
        ri_dmac_data_vld <= i_dmac_data_vld;
        ri_smac_data     <= i_smac_data_vld ? i_smac_data : ri_smac_data;
        ri_smac_data_vld <= i_smac_data_vld;
        ri_vlan_id       <= i_smac_data_vld ? i_vlan_id : ri_vlan_id;
    end
end

// DMAC HASH ʹ���߼���ֱ��ʹ��������Ч�źţ�
always @(posedge i_clk) begin
    if (i_rst) begin
        r_dmac_hash_en  <= 1'b0;
    end else begin
        r_dmac_hash_en  <= i_dmac_data_vld;
    end
end

// SMAC HASH ʹ���߼���ֱ��ʹ��������Ч�źţ�
always @(posedge i_clk) begin
    if (i_rst) begin
        r_smac_hash_en  <= 1'b0;
    end else begin
        r_smac_hash_en  <= i_smac_data_vld;
    end
end

// DMAC HASH ��Ч
always @(posedge i_clk) begin
    if (i_rst) begin
        r_dmac_hash_vld <= 1'b0;
    end else begin
        r_dmac_hash_vld <= r_dmac_hash_en;
    end
end

// SMAC HASH ��Ч
always @(posedge i_clk) begin
    if (i_rst) begin
        r_smac_hash_vld <= 1'b0;
    end else begin
        r_smac_hash_vld <= r_smac_hash_en;
    end
end

always@(posedge i_clk or posedge i_rst ) begin
    if(i_rst) begin
        r_hash_cacl_rst <= 1'd1;
    end else begin
        r_hash_cacl_rst <= r_smac_hash_vld ? 1'd1 : 1'd0;
    end


end

// VLAN ID �����ʹ�ô��ĺ��VLAN ID��
always @(posedge i_clk) begin
    if (i_rst) begin
        ro_vlan_id  <= 12'd0;
    end else begin
        ro_vlan_id  <= r_smac_hash_en ? ri_vlan_id : ro_vlan_id;
    end
end

// DMAC �����ֱ��������ĺ��DMAC��
always @(posedge i_clk) begin
    if (i_rst) begin
        ro_dmac     <= 48'd0;
    end else begin
        ro_dmac     <= r_dmac_hash_en ? ri_dmac_data : ro_dmac;
    end
end

// // DMAC ��Ч���
// always @(posedge i_clk) begin
//     if (i_rst) begin
//         ro_dmac_vld <= 1'b0;
//     end else begin
//         ro_dmac_vld <= r_dmac_hash_vld;
//     end
// end

// DMAC HASH KEY ���
always @(posedge i_clk) begin
    if (i_rst) begin
        ro_dmac_hash_key <= 15'd0;
    end else begin
        ro_dmac_hash_key <= w_dmac_crc_out;
    end
end

// SMAC �����ֱ��������ĺ��SMAC��
always @(posedge i_clk) begin
    if (i_rst) begin
        ro_smac     <= 48'd0;
    end else begin
        ro_smac     <= r_smac_hash_en ? ri_smac_data : ro_smac;
    end
end

// // SMAC ��Ч���
// always @(posedge i_clk) begin
//     if (i_rst) begin
//         ro_smac_vld <= 1'b0;
//     end else begin
//         ro_smac_vld <= r_smac_hash_vld;
//     end
// end

// SMAC HASH KEY ���
always @(posedge i_clk) begin
    if (i_rst) begin
        ro_smac_hash_key <= 15'd0;
    end else begin
        ro_smac_hash_key <= w_smac_crc_out;
    end
end

//---------- HASH ����ģ��ʵ���� ----------
// DMAC HASH���㣺ʹ�ô��ĺ��DMAC��VLAN ID
hash_cacl hash_cacl_u1 (
    .i_data_in      ({i_dmac_data, i_vlan_id}  ),
    .i_crc_en       (i_dmac_data_vld           ),
    .o_crc_out      (w_dmac_crc_out            ),
    .i_rst          (r_hash_cacl_rst           ),
    .i_clk          (i_clk                     )
);

// SMAC HASH���㣺ʹ�ô��ĺ��SMAC��VLAN ID
hash_cacl hash_cacl_u2 (
    .i_data_in      ({i_smac_data, i_vlan_id}  ),
    .i_crc_en       (i_smac_data_vld           ),
    .o_crc_out      (w_smac_crc_out            ),
    .i_rst          (r_hash_cacl_rst           ),
    .i_clk          (i_clk                     )
);

endmodule