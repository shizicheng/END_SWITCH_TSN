`define CPU_MAC
`define MAC1
`define MAC2
`define MAC3
`define MAC4
`define MAC5
`define MAC6
`define MAC7
module swlist#(
    parameter                                                   PORT_NUM                =      8        ,  // �������Ķ˿�??
    parameter                                                   PORT_WIDTH              =      PORT_NUM ,  // �˿�λ�����ڶ˿���
    parameter                                                   PORTBIT_WIDTH           =      clog2(PORT_NUM), // �˿�λ��
    parameter                                                   REG_ADDR_BUS_WIDTH      =      8        ,  // ���� MAC ������üĴ�����??λ��
    parameter                                                   REG_DATA_BUS_WIDTH      =      16       ,  // ���� MAC ������üĴ�������λ??
    parameter                                                   METADATA_WIDTH          =      64       ,  // ��Ϣ����METADATA����λ��
    parameter                                                   PORT_MNG_DATA_WIDTH     =      8        ,  // Mac_port_mng ����λ�� 
    parameter                                                   HASH_DATA_WIDTH         =      15       ,  // ��ϣ�����???��λ��
    parameter                                                   ADDR_WIDTH              =      6        ,  // ��ַ������ 
    parameter                                                   VLAN_ID_WIDTH           =      12       ,  // VLAN IDλ��
    parameter                                                   MAC_ADDR_WIDTH          =      48       ,  // MAC��ַλ��
    parameter                                                   STATIC_RAM_SIZE         =      256      ,  // ��???MAC���λ�� 
    parameter                                                   AGE_SCAN_INTERVAL       =      5        ,  // �ϻ�ɨ��������??
    parameter                                                   SIM_MODE                =      0        ,  // ����ģʽ??1=��???����ģʽ��0=����ģʽ
    parameter                                                   AGE_TIME_WIDTH          =      10       ,
    parameter                                                   CROSS_DATA_WIDTH        =     PORT_MNG_DATA_WIDTH*PORT_NUM // �ۺ�������� 
)(
    input               wire                                    i_clk                               ,   // 250MHz
    input               wire                                    i_rst                               ,   
`ifdef CPU_MAC
    input               wire   [11:0]                           i_vlan_id_cpu                       , // VLAN ID??
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_dmac_cpu_hash_key                 , // Ŀ�� mac �Ĺ�ϣ???
    input               wire   [47 : 0]                         i_dmac_cpu                          , // Ŀ�� mac ��???
    input               wire                                    i_dmac_cpu_vld                      , // dmac_vld
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_smac_cpu_hash_key                 , // ?? mac ��???��Ч��??
    input               wire   [47 : 0]                         i_smac_cpu                          , // ?? mac ��???
    input               wire                                    i_smac_cpu_vld                      , // smac_vld

    output              wire   [PORT_WIDTH - 1:0]               o_tx_cpu_port                       ,
    output              wire                                    o_tx_cpu_port_vld                   ,
    output              wire   [1:0]                            o_tx_cpu_port_broadcast             , // 01:�鲥 10����?? 11:����
`endif
`ifdef MAC1
    input               wire   [11:0]                           i_vlan_id1                          , // VLAN ID??
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_dmac1_hash_key                    , // Ŀ�� mac �Ĺ�ϣ???
    input               wire   [47 : 0]                         i_dmac1                             , // Ŀ�� mac ��???
    input               wire                                    i_dmac1_vld                         , // dmac_vld
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_smac1_hash_key                    , // ?? mac ��???��Ч��??
    input               wire   [47 : 0]                         i_smac1                             , // ?? mac ��???
    input               wire                                    i_smac1_vld                         , // smac_vld

    output              wire   [PORT_WIDTH - 1:0]               o_tx_1_port                         ,
    output              wire                                    o_tx_1_port_vld                     ,
    output              wire   [1:0]                            o_tx_1_port_broadcast               , // 01:�鲥 10����?? 11:����
`endif  
`ifdef MAC2
    input               wire   [11:0]                           i_vlan_id2                          , // VLAN ID??
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_dmac2_hash_key                    , // Ŀ�� mac �Ĺ�ϣ???
    input               wire   [47 : 0]                         i_dmac2                             , // Ŀ�� mac ��???
    input               wire                                    i_dmac2_vld                         , // dmac_vld
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_smac2_hash_key                    , // ?? mac ��???��Ч��??
    input               wire   [47 : 0]                         i_smac2                             , // ?? mac ��???
    input               wire                                    i_smac2_vld                         , // smac_vld

    output              wire   [PORT_WIDTH - 1:0]               o_tx_2_port                         ,
    output              wire                                    o_tx_2_port_vld                     ,
    output              wire   [1:0]                            o_tx_2_port_broadcast               , // 01:�鲥 10����?? 11:����
`endif
`ifdef MAC3
    input               wire   [11:0]                           i_vlan_id3                          , // VLAN ID??
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_dmac3_hash_key                    , // Ŀ�� mac �Ĺ�ϣ???
    input               wire   [47 : 0]                         i_dmac3                             , // Ŀ�� mac ��???
    input               wire                                    i_dmac3_vld                         , // dmac_vld
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_smac3_hash_key                    , // ?? mac ��???��Ч��??
    input               wire   [47 : 0]                         i_smac3                             , // ?? mac ��???
    input               wire                                    i_smac3_vld                         , // smac_vld

    output              wire   [PORT_WIDTH - 1:0]               o_tx_3_port                          ,
    output              wire                                    o_tx_3_port_vld                      ,
    output              wire   [1:0]                            o_tx_3_port_broadcast               , // 01:�鲥 10����?? 11:����
`endif
`ifdef MAC4
    input               wire   [11:0]                           i_vlan_id4                          , // VLAN ID??
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_dmac4_hash_key                    , // Ŀ�� mac �Ĺ�ϣ???
    input               wire   [47 : 0]                         i_dmac4                             , // Ŀ�� mac ��???
    input               wire                                    i_dmac4_vld                         , // dmac_vld
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_smac4_hash_key                    , // ?? mac ��???��Ч��??
    input               wire   [47 : 0]                         i_smac4                             , // ?? mac ��???
    input               wire                                    i_smac4_vld                         , // smac_vld

    output              wire   [PORT_WIDTH - 1:0]               o_tx_4_port                         ,
    output              wire                                    o_tx_4_port_vld                     ,
    output              wire   [1:0]                            o_tx_4_port_broadcast               , // 01:�鲥 10����?? 11:����
`endif
`ifdef MAC5
    input               wire   [11:0]                           i_vlan_id5                          , // VLAN ID??
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_dmac5_hash_key                    , // Ŀ�� mac �Ĺ�ϣ???
    input               wire   [47 : 0]                         i_dmac5                             , // Ŀ�� mac ��???
    input               wire                                    i_dmac5_vld                         , // dmac_vld
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_smac5_hash_key                    , // ?? mac ��???��Ч��??
    input               wire   [47 : 0]                         i_smac5                             , // ?? mac ��???
    input               wire                                    i_smac5_vld                         , // smac_vld

    output              wire   [PORT_WIDTH - 1:0]               o_tx_5_port                         ,
    output              wire                                    o_tx_5_port_vld                     ,
    output              wire   [1:0]                            o_tx_5_port_broadcast               , // 01:�鲥 10����?? 11:����
`endif
`ifdef MAC6
    input               wire   [11:0]                           i_vlan_id6                          , // VLAN ID??
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_dmac6_hash_key                    , // Ŀ�� mac �Ĺ�ϣ???
    input               wire   [47 : 0]                         i_dmac6                             , // Ŀ�� mac ��???
    input               wire                                    i_dmac6_vld                         , // dmac_vld
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_smac6_hash_key                    , // ?? mac ��???��Ч��??
    input               wire   [47 : 0]                         i_smac6                             , // ?? mac ��???
    input               wire                                    i_smac6_vld                         , // smac_vld

    output              wire   [PORT_WIDTH - 1:0]               o_tx_6_port                         ,
    output              wire                                    o_tx_6_port_vld                     ,
    output              wire   [1:0]                            o_tx_6_port_broadcast               , // 01:�鲥 10����?? 11:����
`endif
`ifdef MAC7
    input               wire   [11:0]                           i_vlan_id7                          , // VLAN ID??
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_dmac7_hash_key                    , // Ŀ�� mac �Ĺ�ϣ???
    input               wire   [47 : 0]                         i_dmac7                             , // Ŀ�� mac ��???
    input               wire                                    i_dmac7_vld                         , // dmac_vld
    input               wire   [HASH_DATA_WIDTH - 1 : 0]        i_smac7_hash_key                    , // ?? mac ��???��Ч��??
    input               wire   [47 : 0]                         i_smac7                             , // ?? mac ��???
    input               wire                                    i_smac7_vld                         , // smac_vld

    output              wire   [PORT_WIDTH - 1:0]               o_tx_7_port                         ,
    output              wire                                    o_tx_7_port_vld                     ,
    output              wire   [1:0]                            o_tx_7_port_broadcast               , // 01:�鲥 10����?? 11:����
`endif 
    /*---------------------------------------- �Ĵ������ý�?? -------------------------------------------*/
    // �Ĵ���������??                     
    input               wire                                    i_refresh_list_pulse                , // ˢ�¼Ĵ����б�״???�Ĵ����Ϳ��ƼĴ���??
    input               wire                                    i_switch_err_cnt_clr                , // ˢ�´������??
    input               wire                                    i_switch_err_cnt_stat               , // ˢ�´���״???�Ĵ���
    // �Ĵ���д���ƽӿ�     
    input               wire                                    i_switch_reg_bus_we                 , // �Ĵ���дʹ��
    input               wire   [REG_ADDR_BUS_WIDTH-1:0]         i_switch_reg_bus_we_addr            , // �Ĵ���д��ַ
    input               wire   [REG_DATA_BUS_WIDTH-1:0]         i_switch_reg_bus_we_din             , // �Ĵ���д����
    input               wire                                    i_switch_reg_bus_we_din_v           , // �Ĵ���д����ʹ��
    // �Ĵ��������ƽӿ�     
    input               wire                                    i_switch_reg_bus_rd                 , // �Ĵ�����ʹ��
    input               wire   [REG_ADDR_BUS_WIDTH-1:0]         i_switch_reg_bus_rd_addr            , // �Ĵ�������ַ
    output              wire   [REG_DATA_BUS_WIDTH-1:0]         o_switch_reg_bus_rd_dout            , // �����Ĵ�����??
    output              wire                                    o_switch_reg_bus_rd_dout_v            // ��������Чʹ??
);

// ����ͷ��??
`include "synth_cmd_define.vh"

/*---------------------------------------- clog2���㺯�� -------------------------------------------*/
function integer clog2;
    input integer value;
    integer temp;
    begin
        temp = value - 1;
        for (clog2 = 0; temp > 0; clog2 = clog2 + 1)
            temp = temp >> 1;
    end
endfunction 

// key_arbitģ��������ٲý����??
    wire   [11 : 0]                         w_vlan_id                           ; // VLAN ID�ź�
    wire   [PORT_WIDTH - 1:0]               w_dmac_port                         ; // �ٲ������DMAC�˿�
    wire   [HASH_DATA_WIDTH - 1 : 0]        w_dmac_hash_key                     ; // Ŀ��MAC�Ĺ�ϣ???
    wire   [47 : 0]                         w_dmac                              ; // Ŀ��MAC��???
    wire                                    w_dmac_vld                          ; // DMAC��Ч�ź�
    wire   [HASH_DATA_WIDTH - 1 : 0]        w_smac_hash_key                     ; // ԴMAC�Ĺ�ϣ???
    wire   [47 : 0]                         w_smac                              ; // ԴMAC��???
    wire                                    w_smac_vld                          ; // SMAC��Ч�ź�
    wire   [PORT_NUM - 1:0]                 w_tx_port                           ; // ??�������??
    wire                                    w_tx_port_vld                       ; // ??������˿���Ч��??
    wire   [1:0]                            w_tx_port_broadcast                 ; // 01:�鲥 10����?? 11:����
     
    // DMAC���д�ӿ���??
    wire   [11 : 0]                         w_dmac_item_vlan_id                 ; // DMAC��VLAN ID
    wire   [HASH_DATA_WIDTH-1:0]            w_dmac_item_dmac_addr               ; // DMAC��ַ����
    wire                                    w_dmac_item_dmac_addr_vld           ; // DMAC��ַ������Ч??
    wire   [47:0]                           w_dmac_item_dmac_in                 ; // DMAC����
    wire   [HASH_DATA_WIDTH-1:0]            w_dmac_item_smac_addr               ; // SMAC��ַ����
    wire                                    w_dmac_item_smac_addr_vld           ; // SMAC��ַ������Ч??
    wire   [47:0]                           w_dmac_item_smac_in                 ; // SMAC����
    wire   [PORT_NUM - 1:0]                 w_dmac_item_mac_rx_port             ; // DMAC����˿�
    
    // CLASH��ͻ���д�ӿ���??
    wire   [11 : 0]                         w_clash_item_vlan_id                ; // CLASH��VLAN ID
    wire   [HASH_DATA_WIDTH-1:0]            w_clash_item_dmac_addr              ; // CLASH DMAC��ַ����
    wire                                    w_clash_item_dmac_addr_vld          ; // CLASH DMAC��ַ������Ч??
    wire   [47:0]                           w_clash_item_dmac_in                ; // CLASH DMAC����
    wire   [HASH_DATA_WIDTH-1:0]            w_clash_item_smac_addr              ; // CLASH SMAC��ַ����
    wire                                    w_clash_item_smac_addr_vld          ; // CLASH SMAC��ַ������Ч??
    wire   [47:0]                           w_clash_item_smac_in                ; // CLASH SMAC����
    wire   [PORT_NUM - 1:0]                 w_clash_item_mac_rx_port            ; // CLASH����˿�

    // ������ź�
    wire   [PORT_NUM-1: 0]                  w_smac_tx_port_rslt                 ; // SMAC������˿�����
    wire                                    w_smac_tx_port_vld                  ; // SMAC�������Ч�ź�

    wire                                    w_dmac_find_out_en                  ; // DMAC�������ʹ��
    wire   [PORT_NUM-1:0]                   w_dmac_find_rslt                    ; // DMAC���ҽ���˿�����
    wire                                    w_dmac_find_out_clash               ; // DMAC���ҳ�ͻ��־

    wire   [PORT_NUM-1:0]                   w_clash_tx_port_rslt                ; // ��ͻ�������˿���??
    wire                                    w_clash_tx_port_vld                 ; // ��ͻ��������Ч��??

    // look_up_mng����ź�
    wire   [47 : 0]                         w_lookup_dmac_out                   ; // ����������DMAC
    wire   [11 : 0]                         w_lookup_vlan_id                    ; // ����������VLAN ID
    wire                                    w_lookup_dmac_vld_out               ; // ����������DMAC��Ч�ź�

    // key_arbit��������˿ڵ���??  
`ifdef CPU_MAC
    wire   [PORT_NUM-1: 0]                   w_tx_cpu_port                       ; // CPU�˿����
    wire                                     w_tx_cpu_port_vld                   ; // CPU�˿������Ч
    wire   [1:0]                             w_tx_cpu_port_broadcast             ; // CPU�˿ڹ㲥�������
`endif
`ifdef MAC1
    wire   [PORT_NUM-1: 0]                   w_tx_1_port                         ; // MAC1�˿����
    wire                                     w_tx_1_port_vld                     ; // MAC1�˿������Ч
    wire   [1:0]                             w_tx_1_port_broadcast               ; // MAC1�˿ڹ㲥�������
`endif
`ifdef MAC2
    wire   [PORT_NUM-1: 0]                   w_tx_2_port                         ; // MAC2�˿����
    wire                                     w_tx_2_port_vld                     ; // MAC2�˿������Ч
    wire   [1:0]                             w_tx_2_port_broadcast               ; // MAC2�˿ڹ㲥�������
`endif
`ifdef MAC3
    wire   [PORT_NUM-1: 0]                   w_tx_3_port                         ; // MAC3�˿����
    wire                                     w_tx_3_port_vld                     ; // MAC3�˿������Ч
    wire   [1:0]                             w_tx_3_port_broadcast               ; // MAC3�˿ڹ㲥�������
`endif
`ifdef MAC4
    wire   [PORT_NUM-1: 0]                   w_tx_4_port                         ; // MAC4�˿����
    wire                                     w_tx_4_port_vld                     ; // MAC4�˿������Ч
    wire   [1:0]                             w_tx_4_port_broadcast               ; // MAC4�˿ڹ㲥�������
`endif
`ifdef MAC5
    wire   [PORT_NUM-1: 0]                   w_tx_5_port                         ; // MAC5�˿����
    wire                                     w_tx_5_port_vld                     ; // MAC5�˿������Ч
    wire   [1:0]                             w_tx_5_port_broadcast               ; // MAC5�˿ڹ㲥�������
`endif
`ifdef MAC6
    wire   [PORT_NUM-1: 0]                   w_tx_6_port                         ; // MAC6�˿����
    wire                                     w_tx_6_port_vld                     ; // MAC6�˿������Ч
    wire   [1:0]                             w_tx_6_port_broadcast               ; // MAC6�˿ڹ㲥�������
`endif
`ifdef MAC7
    wire   [PORT_NUM-1: 0]                   w_tx_7_port                         ; // MAC7�˿����
    wire                                     w_tx_7_port_vld                     ; // MAC7�˿������Ч
    wire   [1:0]                             w_tx_7_port_broadcast               ; // MAC7�˿ڹ㲥�������
`endif

    wire        [HASH_DATA_WIDTH-1:0]           w_mac_table_addr                        ;
    wire        [3:0]                           w_fsm_cur_state                         ;

    wire                                        w_table_clear_req                       ;
    wire        [AGE_TIME_WIDTH-1:0]            w_age_time_threshold                    ;
    wire                                        w_table_rd                              ;
    wire        [11:0]                          w_table_raddr                           ;
    wire        [14:0]                          w_table_full_threshold                  ;
    wire        [31:0]                          w_age_scan_interval                     ;

    wire        [57:0]                          w_dmac_list_dout                        ;
    wire        [15:0]                          w_dmac_list_cnt                         ;
    wire                                        w_dmac_list_full_er_stat                ;
    wire        [15:0]                          w_dmac_list_full_er_cnt                 ;

    wire        [14:0]                          w_table_entry_cnt                       ;
    wire        [15:0]                          w_learn_success_cnt                     ;
    wire        [REG_DATA_BUS_WIDTH-1:0]        w_collision_cnt                         ;
    wire        [REG_DATA_BUS_WIDTH-1:0]        w_port_move_cnt                         ;



    // ���˿������??
`ifdef CPU_MAC
    assign o_tx_cpu_port = w_tx_cpu_port[PORT_NUM-1:0];                          // ����CPU�˿����
    assign o_tx_cpu_port_vld = w_tx_cpu_port_vld;                                // ����CPU�˿���Ч�ź�
    assign o_tx_cpu_port_broadcast = w_tx_cpu_port_broadcast;                    // ����CPU�˿ڹ㲥�����ź�
`endif
`ifdef MAC1
    assign o_tx_1_port = w_tx_1_port[PORT_NUM-1:0];                              // ����MAC1�˿����
    assign o_tx_1_port_vld = w_tx_1_port_vld;                                    // ����MAC1�˿���Ч�ź�
    assign o_tx_1_port_broadcast = w_tx_1_port_broadcast;                        // ����MAC1�˿ڹ㲥�����ź�
`endif
`ifdef MAC2
    assign o_tx_2_port = w_tx_2_port[PORT_NUM-1:0];                              // ����MAC2�˿����
    assign o_tx_2_port_vld = w_tx_2_port_vld;                                    // ����MAC2�˿���Ч�ź�
    assign o_tx_2_port_broadcast = w_tx_2_port_broadcast;                        // ����MAC2�˿ڹ㲥�����ź�
`endif
`ifdef MAC3
    assign o_tx_3_port = w_tx_3_port[PORT_NUM-1:0];                              // ����MAC3�˿����
    assign o_tx_3_port_vld = w_tx_3_port_vld;                                    // ����MAC3�˿���Ч�ź�
    assign o_tx_3_port_broadcast = w_tx_3_port_broadcast;                        // ����MAC3�˿ڹ㲥�����ź�
`endif
`ifdef MAC4
    assign o_tx_4_port = w_tx_4_port[PORT_NUM-1:0];                              // ����MAC4�˿����
    assign o_tx_4_port_vld = w_tx_4_port_vld;                                    // ����MAC4�˿���Ч�ź�
    assign o_tx_4_port_broadcast = w_tx_4_port_broadcast;                        // ����MAC4�˿ڹ㲥�����ź�
`endif
`ifdef MAC5
    assign o_tx_5_port = w_tx_5_port[PORT_NUM-1:0];                              // ����MAC5�˿����
    assign o_tx_5_port_vld = w_tx_5_port_vld;                                    // ����MAC5�˿���Ч�ź�
    assign o_tx_5_port_broadcast = w_tx_5_port_broadcast;                        // ����MAC5�˿ڹ㲥�����ź�
`endif
`ifdef MAC6
    assign o_tx_6_port = w_tx_6_port[PORT_NUM-1:0];                              // ����MAC6�˿����
    assign o_tx_6_port_vld = w_tx_6_port_vld;                                    // ����MAC6�˿���Ч�ź�
    assign o_tx_6_port_broadcast = w_tx_6_port_broadcast;                        // ����MAC6�˿ڹ㲥�����ź�
`endif
`ifdef MAC7
    assign o_tx_7_port = w_tx_7_port[PORT_NUM-1:0];                              // ����MAC7�˿����
    assign o_tx_7_port_vld = w_tx_7_port_vld;                                    // ����MAC7�˿���Ч�ź�
    assign o_tx_7_port_broadcast = w_tx_7_port_broadcast;                        // ����MAC7�˿ڹ㲥�����ź�
`endif
    

// �ⲿ����??Ҫ������Ϣ   
key_arbit #(
    .PORT_NUM                   (PORT_NUM                   ),
    .REG_ADDR_BUS_WIDTH         (REG_ADDR_BUS_WIDTH         ),
    .REG_DATA_BUS_WIDTH         (REG_DATA_BUS_WIDTH         ),
    .METADATA_WIDTH             (METADATA_WIDTH             ),
    .PORT_MNG_DATA_WIDTH        (PORT_MNG_DATA_WIDTH        ),
    .HASH_DATA_WIDTH            (HASH_DATA_WIDTH            ) 
) key_arbit_inst (
    .i_clk                      (i_clk                      ),
    .i_rst                      (i_rst                      ),
`ifdef CPU_MAC
    .i_vlan_id_cpu              (i_vlan_id_cpu              ),
    .i_dmac_cpu_hash_key        (i_dmac_cpu_hash_key        ),
    .i_dmac_cpu                 (i_dmac_cpu                 ),
    .i_dmac_cpu_vld             (i_dmac_cpu_vld             ),
    .i_smac_cpu_hash_key        (i_smac_cpu_hash_key        ),
    .i_smac_cpu                 (i_smac_cpu                 ),
    .i_smac_cpu_vld             (i_smac_cpu_vld             ),
    .o_tx_cpu_port              (w_tx_cpu_port              ), 
    .o_tx_cpu_port_vld          (w_tx_cpu_port_vld          ), 
    .o_tx_cpu_port_broadcast    (w_tx_cpu_port_broadcast    ),
`endif
`ifdef MAC1
    .i_vlan_id1                 (i_vlan_id1                 ),
    .i_dmac1_hash_key           (i_dmac1_hash_key           ),
    .i_dmac1                    (i_dmac1                    ),
    .i_dmac1_vld                (i_dmac1_vld                ),
    .i_smac1_hash_key           (i_smac1_hash_key           ),
    .i_smac1                    (i_smac1                    ),
    .i_smac1_vld                (i_smac1_vld                ),
    .o_tx_1_port                (w_tx_1_port                ), 
    .o_tx_1_port_vld            (w_tx_1_port_vld            ), 
    .o_tx_1_port_broadcast      (w_tx_1_port_broadcast      ),
`endif
`ifdef MAC2
    .i_vlan_id2                 (i_vlan_id2                 ),
    .i_dmac2_hash_key           (i_dmac2_hash_key           ),
    .i_dmac2                    (i_dmac2                    ),
    .i_dmac2_vld                (i_dmac2_vld                ),
    .i_smac2_hash_key           (i_smac2_hash_key           ),
    .i_smac2                    (i_smac2                    ),
    .i_smac2_vld                (i_smac2_vld                ),
    .o_tx_2_port                (w_tx_2_port                ), 
    .o_tx_2_port_vld            (w_tx_2_port_vld            ), 
    .o_tx_2_port_broadcast      (w_tx_2_port_broadcast      ),
`endif
`ifdef MAC3
    .i_vlan_id3                 (i_vlan_id3                 ),
    .i_dmac3_hash_key           (i_dmac3_hash_key           ),
    .i_dmac3                    (i_dmac3                    ),
    .i_dmac3_vld                (i_dmac3_vld                ),
    .i_smac3_hash_key           (i_smac3_hash_key           ),
    .i_smac3                    (i_smac3                    ),
    .i_smac3_vld                (i_smac3_vld                ),
    .o_tx_3_port                (w_tx_3_port                ), 
    .o_tx_3_port_vld            (w_tx_3_port_vld            ), 
    .o_tx_3_port_broadcast      (w_tx_3_port_broadcast      ),
`endif
`ifdef MAC4
    .i_vlan_id4                 (i_vlan_id4                 ),
    .i_dmac4_hash_key           (i_dmac4_hash_key           ),
    .i_dmac4                    (i_dmac4                    ),
    .i_dmac4_vld                (i_dmac4_vld                ),
    .i_smac4_hash_key           (i_smac4_hash_key           ),
    .i_smac4                    (i_smac4                    ),
    .i_smac4_vld                (i_smac4_vld                ),
    .o_tx_4_port                (w_tx_4_port                ), 
    .o_tx_4_port_vld            (w_tx_4_port_vld            ), 
    .o_tx_4_port_broadcast      (w_tx_4_port_broadcast      ),
`endif
`ifdef MAC5
    .i_vlan_id5                 (i_vlan_id5                 ),
    .i_dmac5_hash_key           (i_dmac5_hash_key           ),
    .i_dmac5                    (i_dmac5                    ),
    .i_dmac5_vld                (i_dmac5_vld                ),
    .i_smac5_hash_key           (i_smac5_hash_key           ),
    .i_smac5                    (i_smac5                    ),
    .i_smac5_vld                (i_smac5_vld                ),
    .o_tx_5_port                (w_tx_5_port                ), 
    .o_tx_5_port_vld            (w_tx_5_port_vld            ), 
    .o_tx_5_port_broadcast      (w_tx_5_port_broadcast      ),
`endif
`ifdef MAC6
    .i_vlan_id6                 (i_vlan_id6                 ),
    .i_dmac6_hash_key           (i_dmac6_hash_key           ),
    .i_dmac6                    (i_dmac6                    ),
    .i_dmac6_vld                (i_dmac6_vld                ),
    .i_smac6_hash_key           (i_smac6_hash_key           ),
    .i_smac6                    (i_smac6                    ),
    .i_smac6_vld                (i_smac6_vld                ),
    .o_tx_6_port                (w_tx_6_port                ), 
    .o_tx_6_port_vld            (w_tx_6_port_vld            ), 
    .o_tx_6_port_broadcast      (w_tx_6_port_broadcast      ),
`endif
`ifdef MAC7
    .i_vlan_id7                 (i_vlan_id7                 ),
    .i_dmac7_hash_key           (i_dmac7_hash_key           ),
    .i_dmac7                    (i_dmac7                    ),
    .i_dmac7_vld                (i_dmac7_vld                ),
    .i_smac7_hash_key           (i_smac7_hash_key           ),
    .i_smac7                    (i_smac7                    ),
    .i_smac7_vld                (i_smac7_vld                ),
    .o_tx_7_port                (w_tx_7_port                ), 
    .o_tx_7_port_vld            (w_tx_7_port_vld            ), 
    .o_tx_7_port_broadcast      (w_tx_7_port_broadcast      ),
`endif
    // �ٲ����
    .o_dmac_port                (w_dmac_port                ),
    .o_vlan_id                  (w_vlan_id                  ),
    .o_dmac_hash_key            (w_dmac_hash_key            ),
    .o_dmac                     (w_dmac                     ),
    .o_dmac_vld                 (w_dmac_vld                 ),
    .o_smac_hash_key            (w_smac_hash_key            ),
    .o_smac                     (w_smac                     ),
    .o_smac_vld                 (w_smac_vld                 ),
    // ���������
    .i_tx_port                  (w_tx_port                  ),
    .i_tx_port_vld              (w_tx_port_vld              ),
    .i_tx_port_broadcast        (w_tx_port_broadcast        )
);

// ���ٲ�ģ�����룬ͨ����������ַ����������ģ�飬�������ģ�鷵�ز�����������ٲõõ����յĲ���������ظ���һ??
look_up_mng #(
    .HASH_DATA_WIDTH            (HASH_DATA_WIDTH              ),
    .PORT_NUM                   (PORT_NUM                     ),
    .ADDR_WIDTH                 (ADDR_WIDTH                   ),
    .LOCAL_MAC                  (48'h000000000001             )
) look_up_mng_inst (    
    .i_clk                      (i_clk                        ),
    .i_rst                      (i_rst                        ),
    /*------------------------------- KEY�ٲý������ --------------------*/
    .i_vlan_id                  (w_vlan_id                    ), 
    .i_dmac_port                (w_dmac_port                  ),
    .i_dmac_hash_key            (w_dmac_hash_key              ),
    .i_dmac                     (w_dmac                       ),
    .i_dmac_vld                 (w_dmac_vld                   ),
    .i_smac_hash_key            (w_smac_hash_key              ),
    .i_smac                     (w_smac                       ),
    .i_smac_vld                 (w_smac_vld                   ),
    
    .o_tx_port                  (w_tx_port                    ), 
    .o_tx_port_vld              (w_tx_port_vld                ), 
    .o_tx_port_broadcast        (w_tx_port_broadcast          ),
    /*----------------------------- SMAC ���д��?? ------------------------*/         
    .o_dmac                     (w_lookup_dmac_out            ), 
    .o_vlan_id                  (w_lookup_vlan_id             ),
    .o_dmac_vld                 (w_lookup_dmac_vld_out        ), 
    /*----------------------------- DMAC ���д��?? ------------------------*/
    .o_dmac_item_vlan_id        (w_dmac_item_vlan_id          ),
    .o_dmac_item_dmac_addr      (w_dmac_item_dmac_addr        ), 
    .o_dmac_item_dmac_addr_vld  (w_dmac_item_dmac_addr_vld    ), 
    .o_dmac_item_dmac           (w_dmac_item_dmac_in          ), 
    .o_dmac_item_smac_addr      (w_dmac_item_smac_addr        ), 
    .o_dmac_item_smac_addr_vld  (w_dmac_item_smac_addr_vld    ), 
    .o_dmac_item_smac           (w_dmac_item_smac_in          ), 
    .o_dmac_item_mac_rx_port    (w_dmac_item_mac_rx_port      ), 
    /*----------------------------- ��ϣ��ͻ���д��?? -----------------------*/
    .o_clash_item_vlan_id       (w_clash_item_vlan_id         ),
    .o_clash_item_dmac_addr     (w_clash_item_dmac_addr       ), 
    .o_clash_item_dmac_addr_vld (w_clash_item_dmac_addr_vld   ), 
    .o_clash_item_dmac          (w_clash_item_dmac_in         ), 
    .o_clash_item_smac_addr     (w_clash_item_smac_addr       ), 
    .o_clash_item_smac_addr_vld (w_clash_item_smac_addr_vld   ), 
    .o_clash_item_smac          (w_clash_item_smac_in         ), 
    .o_clash_item_mac_rx_port   (w_clash_item_mac_rx_port     ), 
    /*----------------------------- ���Ľ�?? ------------------------------*/
    .i_smac_tx_port_rslt        (w_smac_tx_port_rslt          ), 
    .i_smac_tx_port_vld         (w_smac_tx_port_vld           ), 

    .i_dmac_tx_port_rslt        (w_dmac_find_rslt             ), 
    .i_dmac_lookup_vld          (w_dmac_find_out_en           ), 
    .i_dmac_lookup_clash        (w_dmac_find_out_clash        ), 
	.i_dmac_list_dout           (w_dmac_list_dout             ),  // DMAC�������?? //modify at 12.02

    .i_clash_tx_port_rslt       (w_clash_tx_port_rslt         ), 
    .i_clash_tx_port_vld        (w_clash_tx_port_vld          )  
);

// ��???MAC��������ѧϰMAC��֧���ϻ�����
dmac_mng #(
    .PORT_NUM                   (PORT_NUM                   ),
    .HASH_DATA_WIDTH            (HASH_DATA_WIDTH            ),
    .REG_ADDR_BUS_WIDTH         (REG_ADDR_BUS_WIDTH         ),
    .REG_DATA_BUS_WIDTH         (REG_DATA_BUS_WIDTH         ), 
    .AGE_SCAN_INTERVAL          (AGE_SCAN_INTERVAL          ),
    .SIM_MODE                   (SIM_MODE                   )
) dmac_mng_inst (
    .i_clk                      (i_clk                      ),
    .i_rst                      (i_rst                      ),
    // reg write
    //.i_reg_bus_we               (i_switch_reg_bus_we        ), 
    //.i_reg_bus_addr             (i_switch_reg_bus_we_addr   ), 
    //.i_reg_bus_data             (i_switch_reg_bus_we_din    ), 
    //.i_reg_bus_data_vld         (i_switch_reg_bus_we_din_v  ),
    // reg read
    //.i_reg_bus_re               (i_switch_reg_bus_rd        ), 
    //.i_reg_bus_raddr            (i_switch_reg_bus_rd_addr   ), 
    //.o_reg_bus_rdata            (o_switch_reg_bus_rd_dout   ), 
    //.o_reg_bus_rdata_vld        (o_switch_reg_bus_rd_dout_v ),
    // DMAC/SMAC lookup
    .i_vlan_id                  (w_dmac_item_vlan_id        ), 
    .i_dmac                     (w_dmac_item_dmac_in        ),   
    .i_dmac_hash_addr           (w_dmac_item_dmac_addr      ),   
    .i_dmac_hash_vld            (w_dmac_item_dmac_addr_vld  ),   
    .i_smac                     (w_dmac_item_smac_in        ),   
    .i_smac_hash_addr           (w_dmac_item_smac_addr      ),  
    .i_smac_hash_vld            (w_dmac_item_smac_addr_vld  ),   
    .i_rx_port                  (w_dmac_item_mac_rx_port    ),   
    // lookup output
    .o_dmac_lookup_vld          (w_dmac_find_out_en         ),              
    .o_dmac_tx_port             (w_dmac_find_rslt           ),            
    .o_dmac_lookup_hit          (                           ),         
    .o_lookup_clash             (w_dmac_find_out_clash      ), 
    .o_table_full               (                           ),
    // �Ĵ�??
    .i_table_clear_req          (w_table_clear_req          ),
    .i_age_time_threshold       (w_age_time_threshold       ),
    .i_table_rd                 (w_table_rd                 ),
    .i_table_raddr              (w_table_raddr              ),
    .i_table_full_threshold     (w_table_full_threshold     ),
    .i_age_scan_interval        (w_age_scan_interval        ),
    .o_mac_table_addr           (w_mac_table_addr           ),
    .o_fsm_cur_state            (w_fsm_cur_state            ),
    .o_dmac_list_dout           (w_dmac_list_dout           ),
    .o_dmac_list_cnt            (w_dmac_list_cnt            ),
    .o_dmac_list_full_er_stat   (w_dmac_list_full_er_stat   ),
    .o_dmac_list_full_er_cnt    (w_dmac_list_full_er_cnt    ),
    .o_table_entry_cnt          (w_table_entry_cnt          ),
    .o_learn_success_cnt        (w_learn_success_cnt        ),
    .o_collision_cnt            (w_collision_cnt            ),
    .o_port_move_cnt            (w_port_move_cnt            )
);

/*---------------------------------------- swlist_regs ģ������ -------------------------------------------*/
swlist_regs #(
    .REG_ADDR_BUS_WIDTH         (REG_ADDR_BUS_WIDTH         ),  // �Ĵ�����??λ��
    .REG_DATA_BUS_WIDTH         (REG_DATA_BUS_WIDTH         ),  // �Ĵ�������λ??
    .AGE_TIME_WIDTH             (AGE_TIME_WIDTH             ),  // �ϻ�ʱ��λ��
    .TABLE_FULL_THRESHOLD       (29491                      ),  // MAC������???
    .AGE_SCAN_INTERVAL          (AGE_SCAN_INTERVAL          ),  // �ϻ�ɨ����
    .SIM_MODE                   (SIM_MODE                   )   // ����ģʽ
) u_swlist_regs (
    .i_clk                      (i_clk                      ),  // 250MHzʱ��
    .i_rst                      (i_rst                      ),  // ��λ�ź�
    // �Ĵ���д���ƽӿ�
    .i_reg_bus_we               (i_switch_reg_bus_we        ),  // �Ĵ���дʹ��
    .i_reg_bus_addr             (i_switch_reg_bus_we_addr   ),  // �Ĵ���д��ַ
    .i_reg_bus_data             (i_switch_reg_bus_we_din    ),  // �Ĵ���д����
    .i_reg_bus_data_vld         (i_switch_reg_bus_we_din_v  ),  // �Ĵ���д������Ч
    // �Ĵ��������ƽӿ�
    .i_reg_bus_re               (i_switch_reg_bus_rd        ),  // �Ĵ�����ʹ��
    .i_reg_bus_raddr            (i_switch_reg_bus_rd_addr   ),  // �Ĵ�������ַ
    .o_reg_bus_rdata            (o_switch_reg_bus_rd_dout   ),  // �Ĵ���������(��ʱ����)
    .o_reg_bus_rdata_vld        (o_switch_reg_bus_rd_dout_v ),  // �Ĵ�����������Ч(��ʱ����)

    // MAC�������??
    .i_mac_table_addr           (w_mac_table_addr           ),  // MAC���??
    .i_fsm_cur_state            (w_fsm_cur_state            ),  // ״???����ǰ״???
    .o_table_clear_req          (w_table_clear_req          ),  // �������??
    .o_age_time_threshold       (w_age_time_threshold       ),  // �ϻ�ʱ����???
    .o_table_rd                 (w_table_rd                 ),  // ���ʹ��
    .o_table_raddr              (w_table_raddr              ),  // �����ַ
    .o_table_full_threshold     (w_table_full_threshold     ),
    .o_age_scan_interval        (w_age_scan_interval        ),
    // MAC��״̬��??
    .i_dmac_list_dout           (w_dmac_list_dout           ),  // DMAC�������??
    .i_dmac_list_cnt            (w_dmac_list_cnt            ),  // DMAC���??
    .i_dmac_list_full_er_stat   (w_dmac_list_full_er_stat   ),  // DMAC��������״???
    .i_dmac_list_full_er_cnt    (w_dmac_list_full_er_cnt    ),  // DMAC�����������
    .i_table_entry_cnt          (w_table_entry_cnt          ),  // MAC�������
    .i_learn_success_cnt        (w_learn_success_cnt        ),  // ѧϰ�ɹ�����
    .i_collision_cnt            (w_collision_cnt            ),  // ��ϣ��ͻ����
    .i_port_move_cnt            (w_port_move_cnt            )   // �˿��ƶ�����
);


// ��???MAC������??
// smac_mng #(
//     .DATA_WIDTH                 (VLAN_ID_WIDTH+MAC_ADDR_WIDTH ),
//     .STATIC_RAM_SIZE            (STATIC_RAM_SIZE              ),
//     .REG_ADDR_BUS_WIDTH         (REG_ADDR_BUS_WIDTH           ),
//     .REG_DATA_BUS_WIDTH         (REG_DATA_BUS_WIDTH           )
// ) smac_mng_inst (    
//     .i_sys_clk                  (i_clk                        ),
//     .i_sys_rst                  (i_rst                        ),
//     
//     // reg port    
//     .i_ram_reg_bus_we           (i_switch_reg_bus_we          ), 
//     .i_ram_reg_bus_we_addr      (i_switch_reg_bus_we_addr     ),
//     .i_ram_reg_bus_we_din       (i_switch_reg_bus_we_din      ),
//     .i_ram_reg_bus_we_din_v     (i_switch_reg_bus_we_din_v    ),
//     
//     .i_ram_reg_bus_rd           (i_switch_reg_bus_rd          ),
//     .i_ram_reg_bus_rd_addr      (i_switch_reg_bus_rd_addr     ),
//     .o_ram_reg_bus_we_din       (o_switch_reg_bus_rd_dout     ),
//     .o_ram_reg_bus_we_din_v     (o_switch_reg_bus_rd_dout_v   ),
//     
//     // input data port    
//     .i_vlan_id                  (w_vlan_id                    ),
//     .i_query_data               (w_lookup_dmac_out            ), 
//     .i_query_valid              (w_lookup_dmac_vld_out        ),
//     
//     // output data port    
//     .o_port_vector              (w_smac_tx_port_rslt          ),
//     .o_port_vector_valid        (w_smac_tx_port_vld           )
// );


// HASH��ͻ?? �����???MAC����ֳ�ͻ�����Գ�ͻ��Ĳ����Ϊ׼ 
// clash_mac_mng #(
//     .DATA_WIDTH                 (VLAN_ID_WIDTH+MAC_ADDR_WIDTH ),
//     .STATIC_RAM_SIZE            (STATIC_RAM_SIZE              ),
//     .REG_ADDR_BUS_WIDTH         (REG_ADDR_BUS_WIDTH           ),
//     .REG_DATA_BUS_WIDTH         (REG_DATA_BUS_WIDTH           )
// ) clash_mac_mng_inst (
//     .i_sys_clk                  (i_clk                        ),
//     .i_sys_rst                  (i_rst                        ),
// 
//     // reg port
//     .i_ram_reg_bus_we           (i_switch_reg_bus_we          ), 
//     .i_ram_reg_bus_we_addr      (i_switch_reg_bus_we_addr     ),
//     .i_ram_reg_bus_we_din       (i_switch_reg_bus_we_din      ),
//     .i_ram_reg_bus_we_din_v     (i_switch_reg_bus_we_din_v    ),
// 
//     .i_ram_reg_bus_rd           (i_switch_reg_bus_rd          ),
//     .i_ram_reg_bus_rd_addr      (i_switch_reg_bus_rd_addr     ),
//     .o_ram_reg_bus_we_din       (o_switch_reg_bus_rd_dout     ),
//     .o_ram_reg_bus_we_din_v     (o_switch_reg_bus_rd_dout_v   ),
// 
//     // input data port
//     .i_query_data               (w_clash_item_dmac_in          ), 
//     .i_query_valid              (w_clash_item_dmac_addr_vld    ),
// 
//     // output data port
//     .o_port_vector              (w_clash_tx_port_rslt          ),
//     .o_port_vector_valid        (w_clash_tx_port_vld           )
// );

endmodule
