module rx_forward_mng#(
    parameter                                                   PORT_NUM                =      4        ,  // �������Ķ˿���
    parameter                                                   PORT_MNG_DATA_WIDTH     =      8        ,  // Mac_port_mng ����λ��
    parameter                                                   METADATA_WIDTH          =      81       ,  // ��Ϣ��λ��
	parameter                                                   PORT_INDEX              =      0        , 
    parameter                                                   CROSS_DATA_WIDTH        =     PORT_MNG_DATA_WIDTH*PORT_NUM // �ۺ��������
)(
    input               wire                                    i_clk                              ,   // 250MHz
    input               wire                                    i_rst                              ,
    /*---------------------------------------- ����ת����صļĴ��� -------------------------------------------*/
    input              wire                                     i_port_rxmac_down_regs             , // �˿ڽ��շ���MAC�ر�ʹ��
    input              wire                                     i_port_broadcast_drop_regs         , // �˿ڹ㲥֡����ʹ��
    input              wire                                     i_port_multicast_drop_regs         , // �˿��鲥֡����ʹ��
    input              wire                                     i_port_loopback_drop_regs          , // �˿ڻ���֡����ʹ��
    input              wire   [47:0]                            i_port_mac_regs                    , // �˿ڵ� MAC ��ַ
    input              wire                                     i_port_mac_vld_regs                , // ʹ�ܶ˿� MAC ��ַ��Ч
    input              wire   [7:0]                             i_port_mtu_regs                    , // MTU����ֵ
    input              wire   [PORT_NUM-1:0]                    i_port_mirror_frwd_regs            , // ����ת���Ĵ���������Ӧ�Ķ˿���1���򱾶˿ڽ��յ����κ�ת������֡������ת��ֵ����1�Ķ˿�
    input              wire   [15:0]                            i_port_flowctrl_cfg_regs           , // ������������                                                                        
    input              wire   [4:0]                             i_port_rx_ultrashortinterval_num   , // ֡���                                                                          
    /*---------------------------------------- rx_frm_info_mng input ����Ϣ�� -------------------------------------------*/
    input              wire                                     i_rtag_flag                        , // rtag��־ -> CB�ı���    
    input              wire   [15:0]                            i_rtag_sequence                    , // [80:65] : CBЭ�� R-TAG�ֶ�
    input              wire   [1:0]                             i_port_speed                       , // [64:63](2bit) : port_speed 
    input              wire   [2:0]                             i_vlan_pri                         , // [62:60](3bit) : vlan_pri 
    input              wire                                     i_frm_vlan_flag                    , // [27](1bit) : frm_vlan_flag
    // input              wire   [PORT_NUM-1:0]                    i_rx_port                          , // [26:19](8bit) : ����˿ڣ�bitmap��ʾ
    input              wire                                     i_frm_discard                      , // crc�Ƿ���ȷ���Ƿ���
    input              wire                                     i_frm_qbu                          , // [11](1bit) : �Ƿ�Ϊ�ؼ�֡(Qbu)
    // // �ڲ���Ϣ����ʹ�ã�����Ϊmetadata�ֶ� 
    // input              wire                                     i_frm_info_vld                     , // ֡��Ϣ��Ч 
    // input              wire                                     i_broadcast_frm_en                 , // �㲥֡ 
    // input              wire                                     i_multicast_frm_en                 , // �鲥֡ 
    // input              wire                                     i_mac_time_irq                      , // ��ʱ����ж��ź�
    // input              wire   [7:0]                             i_mac_frame_seq                     , // ֡���к�
    input              wire   [6:0]                             i_timestamp_addr                   , // ��ʱ����洢�� RAM ��ַ 
    input              wire   [15:0]                            i_ethertype                        , // ��̫�������ֶ�  
    input              wire                                     i_info_valid                       ,
    /*---------------------------------------- ���ģ����ݹ�ϣֵ���صļ����� ----------------------------------*/
    input              wire    [PORT_NUM-1:0]                  i_swlist_tx_port                    , // ���Ͷ˿���Ϣ   
    input              wire   [1:0]                            i_swlist_port_broadcast             , // 01:�鲥 10���㲥 11:����
    input              wire                                    i_swlist_vld                        , // ��Чʹ���ź�                                   
    /*---------------------------------------- ACL ƥ���������ֶ� ------------------------------ -------------*/
    input              wire                                    i_acl_vld                           , // aclƥ������Ч����ź�
    input              wire    [2:0]                           i_acl_action                        , // ACL����: 000-���� 001-���� 010-�ض���
    input              wire                                    i_acl_cb_frm                        , // CBЭ��֡��־
    input              wire    [7:0]                           i_acl_cb_streamhandle               , // stream_handleֵ(8bit)
    input              wire    [2:0]                           i_acl_flow_ctrl                     , // ��������: 00-100% 01-50% 10-25% 11-12.5%
    input              wire    [7:0]                           i_acl_forwardport                   , // ת���˿�bitmap  
    // input              wire                                    i_acl_find_match                   , // �Ƿ�ƥ�䵽��ȷ����Ŀ
    // input              wire   [7:0]                            i_acl_frmtype                      , // ƥ�������֡����
    // input              wire   [15:0]                           i_acl_fetch_info                   , // �������� 
    
    // input              wire   [1:0]                            i_frm_cb_op                         , // [14:13](2bit) :[0]:1��ʾCBҵ��֡��[0]:0��ʾ��CBҵ��֡  [1]��1 �� rtag ��ǩ [1]��0 �� rtag ��ǩ ok   
    // /*---------------------------------------- �� PORT �ۺ����������� -------------------------------------------*/
    // input              wire                                    i_mac_port_link                    , // �˿ڵ�����״̬
    // input              wire   [1:0]                            i_mac_port_speed                   , // �˿�������Ϣ��00-10M��01-100M��10-1000M��10-10G 

    input              wire   [PORT_MNG_DATA_WIDTH-1:0]        i_mac_port_axi_data                 , // �˿������������λ��ʾcrcerr
    input              wire   [15:0]                           i_mac_axi_data_user                 , // �Ƿ�ؼ�֡ + ���ĳ���
    input              wire   [(PORT_MNG_DATA_WIDTH/8)-1:0]    i_mac_axi_data_keep                 , // �˿����������룬��Ч�ֽ�ָʾ
    input              wire                                    i_mac_axi_data_valid                , // �˿�������Ч
    output             wire                                    o_mac_axi_data_ready                , // �������߾ۺϼܹ���ѹ��ˮ���ź�
    input              wire                                    i_mac_axi_data_last                 , // ������������ʶ
    // /*---------------------------------------- �� PORT �ۺ���������� -------------------------------------------*/
    // output             wire                                    o_mac_port_link                    , // �˿ڵ�����״̬
    // output             wire   [1:0]                            o_mac_port_speed                   , // �˿�������Ϣ��00-10M��01-100M��10-1000M��10-10G 
    output             wire   [PORT_MNG_DATA_WIDTH-1:0]        o_mac_port_axi_data                 , // �˿������������λ��ʾcrcerr
    output             wire   [15:0]                           o_mac_axi_data_user                 , // �Ƿ�ؼ�֡ + ���ĳ���
    output             wire   [(PORT_MNG_DATA_WIDTH/8)-1:0]    o_mac_axi_data_keep                 , // �˿����������룬��Ч�ֽ�ָʾ
    output             wire                                    o_mac_axi_data_valid                , // �˿�������Ч
    input              wire                                    i_mac_axi_data_ready                , // �������߾ۺϼܹ���ѹ��ˮ���ź�
    output             wire                                    o_mac_axi_data_last                 , // ������������ʶ
    /*---------------------------------------- �� PORT �ۺ���Ϣ�� -------------------------------------------*/
    output             wire   [METADATA_WIDTH-1:0]             o_cross_metadata                    , // �ۺ����� metadata ����
    output             wire                                    o_cross_metadata_valid              , // �ۺ����� metadata ������Ч�ź�
    output             wire                                    o_cross_metadata_last               , // ��Ϣ��������ʶ
    input              wire                                    i_cross_metadata_ready              , // ����ģ�鷴ѹ��ˮ�� 
    /*---------------------------------------- ��ϼĴ��� -------------------------------------------*/
    output             wire                                    o_port_rx_ultrashort_frm            , // �˿ڽ��ճ���֡(С��64�ֽ�)
    output             wire                                    o_port_rx_overlength_frm            , // �˿ڽ��ճ���֡(����MTU�ֽ�)
    output             wire                                    o_port_rx_crcerr_frm                , // �˿ڽ���CRC����֡
    output             wire  [15:0]                            o_port_rx_loopback_frm_cnt          , // �˿ڽ��ջ���֡������ֵ
    output             wire  [15:0]                            o_port_broadflow_drop_cnt           , // �˿ڽ��յ��㲥������������֡������ֵ
    output             wire  [15:0]                            o_port_multiflow_drop_cnt           , // �˿ڽ��յ��鲥������������֡������ֵ
    output             wire  [15:0]                            o_port_diag_state                     // �˿�״̬�Ĵ�����������Ĵ�����˵������ 
);

   /*
        metadata ������� (��λ��81bit)
            
            [80:65](16bit): CBЭ�� R-TAG�ֶ� ok
            [64:63](2bit) : port_speed ok
            [62:60](3bit) : vlan_pri ok
            [59:52](8bit) : tx_prot (�ں�ACLת���˿�) ok 
            [51:44](8bit) : acl_frmtype ok
            [43:36](8bit) : stream_handle��CBЭ������ʶ ok
            [35:28](8bit) : �����ֶ�
            [27](1bit)    : frm_vlan_flag ok
            [26:19](8bit) : ����˿ڣ�bitmap��ʾ ok
            [18:15](4bit) : ����
            [14:13](2bit) : ��ʶ��ƥ�䣬[1]:rtag_flag [0]:cb_frm ok 
            [12](1bit)    : ����λ(��ACL action����) ok
            [11](1bit)    : �Ƿ�Ϊ�ؼ�֡(Qbu) ok
            [10:4](7bit)  : time_stamp_addr������ʱ����ĵ�ַ��Ϣ ok
            [3:0](4bit)   : ����
    */
/*--------- �ź������� --------*/

// FIFO��ز�������
localparam FIFO_DEPTH       = 30                                                                ;
localparam FIFO_WIDTH       = PORT_MNG_DATA_WIDTH + (PORT_MNG_DATA_WIDTH/8) + 1                ; // data + keep + last
localparam FIFO_CNT_WIDTH   = 5                                                                 ; // log2(30) ����ȡ��

// FIFO����ź�
wire                                    w_fifo_wr_en                    ; // FIFOдʹ��
wire    [FIFO_WIDTH-1:0]                w_fifo_din                      ; // FIFOд������
wire                                    w_fifo_full                     ; // FIFO���ź�
wire                                    w_fifo_rd_en                    ; // FIFO��ʹ��
wire    [FIFO_WIDTH-1:0]                w_fifo_dout                     ; // FIFO��������
wire                                    w_fifo_empty                    ; // FIFO���ź�
wire    [FIFO_CNT_WIDTH-1:0]            w_fifo_data_cnt                 ; // FIFO���ݼ���

// FIFO������ݽ��
wire    [PORT_MNG_DATA_WIDTH-1:0]       w_fifo_out_data                 ; // FIFO���������
wire    [(PORT_MNG_DATA_WIDTH/8)-1:0]   w_fifo_out_keep                 ; // FIFO�����keep
wire                                    w_fifo_out_last                 ; // FIFO�����last

// user�źŻ��棨ÿ֡��һ�ģ�
reg                                     r_fifo_rd_en                    ;
reg     [15:0]                          r_frame_user                    ; // �����user�ź�

// ����ģ�����wire�ź�
wire    [31:0]                          w_recive_package                ; // ���հ�����
wire    [31:0]                          w_recive_package_multi          ; // ���հ���������
wire    [31:0]                          w_send_package                  ; // ���Ͱ�����
wire    [31:0]                          w_send_package_multi            ; // ���Ͱ���������
wire    [PORT_MNG_DATA_WIDTH-1:0]       w_flow_data_out                 ; // ���غ��������
wire    [(PORT_MNG_DATA_WIDTH/8)-1:0]   w_flow_data_keep_out            ; // ���غ���������
wire                                    w_flow_valid_out                ; // ���غ�������Ч
wire                                    w_flow_ready                 ; // ����ģ��ready
wire                                    w_flow_last_out                 ; // ���غ�last�ź�

// ����ģ������ѡ���ź�
wire    [PORT_MNG_DATA_WIDTH-1:0]       w_flow_ctrl_input_data          ; // ����ģ����������ѡ��
wire    [(PORT_MNG_DATA_WIDTH/8)-1:0]   w_flow_ctrl_input_keep          ; // ����ģ����������ѡ��
wire                                    w_flow_ctrl_input_valid         ; // ����ģ��������Чѡ��
wire                                    w_flow_ctrl_input_last          ; // ����ģ������lastѡ��

// �����ж����������ź�
reg                                     r_acl_match_flow_type           ; // ACLƥ������֡����
reg                                     r_flow_ctrl_enable              ; // ������ʹ��

// ���������ź�
reg     [2:0]                           ri_flow_ctrl_select             ; // �������ô���

// ֡�����ж�����߼�
wire    [7:0]                           w_frm_type                      ; // ������̫�������жϵ�֡����

//-------------------- ���������� --------------------
// �����źŴ��� 
reg                                     ri_mac_axi_data_valid           ;
reg     [PORT_MNG_DATA_WIDTH-1:0]       ri_mac_port_axi_data            ;
reg     [(PORT_MNG_DATA_WIDTH/8)-1:0]   ri_mac_axi_data_keep            ;
reg                                     ri_mac_axi_data_last            ;
reg     [15:0]                          ri_mac_axi_data_user            ;
reg     [15:0]                          ri_rtag_sequence                ;
reg                                     ri_frm_vlan_flag                ;
reg     [2:0]                           ri_vlan_pri                     ;
reg     [PORT_NUM-1:0]                  r_rx_port                       ;
reg     [7:0]                           ri_acl_frmtype                  ;
reg                                     ri_acl_vld                      ; 
// reg     [15:0]                          ri_acl_fetch_info               ;
reg     [1:0]                           ri_frm_cb_op                    ;
reg                                     ri_frm_qbu                      ;
reg     [6:0]                           ri_timestamp_addr               ;
reg     [1:0]                           ri_port_speed                   ;
reg     [15:0]                          ri_ethertype                    ; // ��̫�����ʹ���
reg     [PORT_NUM-1:0]                  ri_swlist_tx_port               ;
reg                                     ri_swlist_vld                   ;
reg                                     ri_frm_discard                  ;
reg     [7:0]                           ri_tx_prot                      ; // metadata�����ֶ�
reg     [3:0]                           ri_qos_policy                   ; // metadata�����ֶ�
reg                                     ri_discard                      ; // metadata����λ
reg     [15:0]                          ri_port_flowctrl_cfg_regs       ; // �������üĴ�������
reg     [2:0]                           ri_acl_action                   ; // ACL�������ʹ���
reg                                     ri_acl_cb_frm                   ; // ACL CBЭ��֡��־����
reg                                     ri_rtag_flag                    ; // RTAG��־����
reg     [7:0]                           ri_acl_cb_streamhandle          ; // ACL stream_handle����
reg     [1:0]                           ri_acl_flow_ctrl                ; // ACL�������ô���
reg     [7:0]                           ri_acl_forwardport              ; // ACLת���˿ڴ���

// ���ش������
reg                                     r_need_flow_ctrl                ;
reg                                     r_need_flow_ctrl_d1             ;

// metadata���
reg     [METADATA_WIDTH-1:0]            ro_cross_metadata               ;
reg                                     ro_cross_metadata_valid         ;
reg                                     ro_cross_metadata_last          ;

// ���������
reg     [PORT_MNG_DATA_WIDTH-1:0]       ro_mac_port_axi_data            ;
reg     [(PORT_MNG_DATA_WIDTH/8)-1:0]   ro_mac_axi_data_keep            ;
reg                                     ro_mac_axi_data_valid           ;
reg                                     ro_mac_axi_data_last            ;
reg     [15:0]                          ro_mac_axi_data_user            ;

// metadata_valid���Ʊ�־λ
reg                                     r_swlist_vld_flag               ; // swlist_vld������־
reg                                     r_acl_vld_flag                  ; // acl_vld������־
wire                                    w_both_vld_ready                ; // ����vld���Ѵ���
wire                                    w_discard                       ;

// FIFO��ȡ����
reg                                     r_lookup_done                   ; // �����ɱ�־
reg                                     r_frame_start                   ; // ֡��ʼ��־
always @(posedge i_clk) begin
    if (i_rst) begin
        ri_mac_axi_data_valid   <= 1'b0;
        ri_mac_port_axi_data    <= {PORT_MNG_DATA_WIDTH{1'b0}};
        ri_mac_axi_data_keep    <= {(PORT_MNG_DATA_WIDTH/8){1'b0}};
        ri_mac_axi_data_last    <= 1'b0;
        ri_mac_axi_data_user    <= 16'd0;
        ri_rtag_sequence        <= 16'd0;
        ri_frm_vlan_flag        <= 1'b0;
        ri_vlan_pri             <= 3'd0;
        ri_acl_frmtype          <= 8'd0;
        ri_acl_vld              <= 1'b0; 
        ri_frm_cb_op            <= 2'd0;
        ri_frm_qbu              <= 1'b0;
        ri_timestamp_addr       <= 8'd0;
        ri_port_speed           <= 2'd0;
        ri_ethertype            <= 16'd0;
        ri_swlist_tx_port       <= {PORT_NUM{1'b0}};
        ri_swlist_vld           <= 1'b0;
        ri_frm_discard          <= 1'b0;
        ri_tx_prot              <= 8'd0;
        ri_qos_policy           <= 4'd0;
        ri_discard              <= 1'b0;
        ri_port_flowctrl_cfg_regs <= 16'd0;
        ri_acl_action           <= 3'd0;
        ri_acl_cb_frm           <= 1'b0;
        ri_rtag_flag            <= 1'b0;
        ri_acl_cb_streamhandle  <= 8'd0;
        ri_acl_flow_ctrl        <= 2'd0;
        ri_acl_forwardport      <= 8'd0; 
    end else begin
        ri_mac_axi_data_valid   <= i_mac_axi_data_valid;
        ri_mac_port_axi_data    <= i_mac_port_axi_data;
        ri_mac_axi_data_keep    <= i_mac_axi_data_keep;
        ri_mac_axi_data_last    <= i_mac_axi_data_last;
        ri_mac_axi_data_user    <= i_mac_axi_data_user;
        ri_rtag_flag            <= i_rtag_flag == 1'd1 || (ri_rtag_flag == 1'd1 && i_mac_axi_data_valid == 1'd1) ? 1'd1 : 1'd0;//ri_mac_axi_data_last ? 1'd0 : ri_rtag_flag
        ri_rtag_sequence        <= i_info_valid ? i_rtag_sequence : ri_rtag_sequence;
        ri_frm_vlan_flag        <= i_info_valid ? i_frm_vlan_flag : ri_frm_vlan_flag;
        ri_vlan_pri             <= i_info_valid ? i_vlan_pri      : ri_vlan_pri     ;
        ri_acl_frmtype          <= w_frm_type;
        ri_acl_vld              <= i_acl_vld; 
        ri_frm_cb_op            <= {ri_rtag_flag, ri_acl_cb_frm}; // [1]:rtag_flag [0]:cb_frm
        ri_frm_qbu              <= i_info_valid ? i_frm_qbu : ri_frm_qbu;
        ri_timestamp_addr       <= i_info_valid ? i_timestamp_addr : ri_timestamp_addr;
        ri_port_speed           <= i_info_valid ? i_port_speed : ri_port_speed;
        ri_ethertype            <= i_info_valid ? i_ethertype  : ri_ethertype ;
        ri_swlist_tx_port       <= i_swlist_vld ? i_swlist_tx_port : ri_swlist_tx_port; // ACLת���˿�����
        ri_swlist_vld           <= i_swlist_vld;
        ri_frm_discard          <= i_info_valid ? i_frm_discard : ri_frm_discard;
        ri_tx_prot              <= (ri_acl_forwardport != 8'd0) ? ri_acl_forwardport[PORT_NUM-1:0] : ri_swlist_tx_port; // ACLת���˿�����  
        ri_qos_policy           <= 4'd1;  
        ri_discard              <= i_info_valid ? i_frm_discard : ri_discard;
        // ri_discard              <= (ri_acl_action == 3'b001) ? 1'b1 : i_frm_discard; // ACL action=001Ϊ����
        ri_port_flowctrl_cfg_regs <= i_port_flowctrl_cfg_regs       ;
        ri_acl_action           <= i_acl_vld ? i_acl_action          : ri_acl_action          ;
        ri_acl_cb_frm           <= i_acl_vld ? i_acl_cb_frm          : ri_acl_cb_frm          ;
        ri_acl_cb_streamhandle  <= i_acl_vld ? i_acl_cb_streamhandle : ri_acl_cb_streamhandle ;
        ri_acl_flow_ctrl        <= i_acl_vld ? i_acl_flow_ctrl       : ri_acl_flow_ctrl       ;
        ri_acl_forwardport      <= i_acl_vld ? i_acl_forwardport     : ri_acl_forwardport     ; 
    end
end

assign w_discard = (ri_acl_action == 3'b001) ? 1'b1 : ri_discard;

// ���ն˿ڱ�ʶ�����ڲ���PORT_INDEX��
always @(posedge i_clk) begin
    if (i_rst) begin
        r_rx_port <= {PORT_NUM{1'b0}};
    end else begin
        r_rx_port <= 1'b1 << PORT_INDEX[2:0];
    end
end
 
//-------------------- ֡�����ж�����߼� --------------------
// ������̫�������ж�֡����
// 0x88F7: 802.1AS (PTP) -> frm_type = 1
// 0x88CC: LLDP          -> frm_type = 2  
// 0x010B: RSTP          -> frm_type = 3
// ����:                 -> frm_type = 0
assign w_frm_type = (i_ethertype == 16'h88F7) ? 8'd1 :
                    (i_ethertype == 16'h88CC) ? 8'd2 :
                    (i_ethertype == 16'h010B) ? 8'd3 : 
                    8'd0;

//-------------------- ���������߼� --------------------
// ��������ƴ�ӣ�ACL�������ȣ����ACL��Ч���������ò�Ϊ0��ʹ��ACL���أ�����ʹ�üĴ�������
// [1:0]: ���صȼ�ѡ�� (00=100%, 01=50%, 10=25%, 11=12.5%)
always @(posedge i_clk) begin
    if (i_rst)
        ri_flow_ctrl_select <= 3'd0;
    else
        ri_flow_ctrl_select <= (i_acl_vld == 1'b1 && i_acl_flow_ctrl != 3'b00) ? i_acl_flow_ctrl : ri_port_flowctrl_cfg_regs[2:0];
end

//-------------------- �����ж��߼� --------------------
// ACLƥ������֡�����ж�
always @(posedge i_clk) begin
    if (i_rst)
        r_acl_match_flow_type <= 1'b0;
    else
        r_acl_match_flow_type <= (ri_acl_vld == 1'b1 && ri_acl_frmtype == 8'h01) ? 1'b1 : 1'b0;
end

// ������ʹ���ж�
always @(posedge i_clk) begin
    if (i_rst)
        r_flow_ctrl_enable <= 1'b0;
    else
        r_flow_ctrl_enable <= 1'd1;  // ���ԣ�r_flow_ctrl_enable <= (ri_port_flowctrl_cfg_regs[12] == 1'b1) ? 1'b1 : 1'b0;
end

// ���ش���ʹ�ܣ�ACLƥ������֡���� && ������ʹ��  // ���ǵ���������
always @(posedge i_clk) begin
    if (i_rst) begin
        r_need_flow_ctrl <= 1'b0;
    end else begin
        // r_need_flow_ctrl <= 1'b0; // ����
        r_need_flow_ctrl <= (i_swlist_port_broadcast != 2'd0 && r_flow_ctrl_enable == 1'b1) ? 1'b1 :
                            (ro_mac_axi_data_last ? 1'b0 : r_need_flow_ctrl); 
    end
end

always @(posedge i_clk) begin
     r_need_flow_ctrl_d1 <=  r_need_flow_ctrl;
end

//-------------------- FIFOд���߼� --------------------
// FIFOд��ʹ�ܣ�����������Ч��FIFOδ��
assign w_fifo_wr_en = i_mac_axi_data_valid && !w_fifo_full;

// FIFOд�����ݴ����data + keep + last (������user)
assign w_fifo_din = {i_mac_axi_data_last, i_mac_axi_data_keep, i_mac_port_axi_data};

//-------------------- user�źŻ����߼� --------------------
// ���֡��ʼ����һ����Ч����ǰ����Ч
always @(posedge i_clk) begin
    if (i_rst)
        r_frame_start <= 1'b0;
    else
        r_frame_start <= (!ri_mac_axi_data_valid && i_mac_axi_data_valid);
end

// ��֡��ʼʱ����user�ź�
always @(posedge i_clk) begin
    if (i_rst)
        r_frame_user <= 16'd0;
    else if (r_frame_start)
        r_frame_user <= {3'b000,ri_acl_cb_frm,i_mac_axi_data_user[11:0]};
end

//-------------------- FIFO��ȡ�߼� --------------------
// �����ɱ�־����i_swlist_vld����ʱ����ʾ������
always @(posedge i_clk) begin
    if (i_rst)
        r_lookup_done <= 1'b0;
    else
        r_lookup_done <= i_swlist_vld ? 1'b1 : (w_fifo_empty ? 1'b0 : r_lookup_done);
end

// FIFO��ȡʹ�ܣ������� && FIFO�ǿ� && ����ready
assign w_fifo_rd_en = r_lookup_done && !w_fifo_empty && 
                      ((r_need_flow_ctrl == 1'b1) ? w_flow_ready : i_mac_axi_data_ready);

// FIFO������ݽ��
assign w_fifo_out_data = w_fifo_dout[PORT_MNG_DATA_WIDTH-1:0];
assign w_fifo_out_keep = w_fifo_dout[PORT_MNG_DATA_WIDTH + (PORT_MNG_DATA_WIDTH/8) - 1 : PORT_MNG_DATA_WIDTH];
assign w_fifo_out_last = w_fifo_dout[FIFO_WIDTH-1];

always @(posedge i_clk) begin  
    r_fifo_rd_en <= w_fifo_rd_en;
end
//-------------------- FIFOģ��ʵ���� --------------------
sync_fifo #(
    .DEPTH                  ( FIFO_DEPTH                )  ,
    .WIDTH                  ( FIFO_WIDTH                )  ,
    .ALMOST_FULL_THRESHOLD  ( 1                         )  ,
    .ALMOST_EMPTY_THRESHOLD ( 1                         )  ,
    .FLOP_DATA_OUT          ( 0                         )  , // ʹ��stdģʽ
    .RAM_STYLE              ( 0                         )    // ʹ��Distributed RAM��С����FIFO��
) u_data_fifo (
    .i_clk                  ( i_clk                     )  ,
    .i_rst                  ( i_rst                     )  ,
    .i_wr_en                ( w_fifo_wr_en              )  ,
    .i_din                  ( w_fifo_din                )  ,
    .o_full                 ( w_fifo_full               )  ,
    .i_rd_en                ( w_fifo_rd_en              )  ,
    .o_dout                 ( w_fifo_dout               )  ,
    .o_empty                ( w_fifo_empty              )  ,
    .o_almost_full          (                           )  , // δʹ��
    .o_almost_empty         (                           )  , // δʹ��
    .o_data_cnt             ( w_fifo_data_cnt           )
);

//-------------------- ����ģ������ѡ���߼� --------------------
// ��FIFO������������������ģ���ֱ�����
assign w_flow_ctrl_input_data  = r_need_flow_ctrl_d1  == 1'd1 && r_fifo_rd_en == 1'd1 ? w_fifo_out_data : {PORT_MNG_DATA_WIDTH{1'b0}};
assign w_flow_ctrl_input_keep  = r_need_flow_ctrl_d1  == 1'd1 && r_fifo_rd_en == 1'd1 ? w_fifo_out_keep : {(PORT_MNG_DATA_WIDTH/8){1'b0}};
assign w_flow_ctrl_input_valid = r_need_flow_ctrl_d1 ? r_fifo_rd_en    : 1'd0;// FIFO��ȡʱ������Ч
assign w_flow_ctrl_input_last  = r_need_flow_ctrl_d1  == 1'd1 && r_fifo_rd_en == 1'd1 ? w_fifo_out_last : 1'd0;

//-------------------- ����ģ��ʵ���� --------------------
// ���ض�֡���������ش���
flow_driver#(
    .SIM_MODE               ( "TRUE"                )  ,
    .REG_DATA_WIDTH         ( 16                    )  ,
    .PORT_MNG_DATA_WIDTH    ( PORT_MNG_DATA_WIDTH   )  ,
    .CLOCK_PERIOD           ( 250_000_000           ) 
) flow_driver_inst (                                       
    .i_sys_clk              ( i_clk                 )  ,
    .i_sys_rst              ( i_rst                 )  ,

    .i_pluse_clk            ( i_clk                 )  , // ʹ��ϵͳʱ��250MHz
    .i_pluse_rst            ( i_rst                 )  ,

    .i_port_rate            ( ri_port_speed         )  , // �˿�����: 00-100M 01-1000M 10-2500M 11-10G
    .i_flow_ctrl_select     (3'd0),//( ri_flow_ctrl_select   )  , // ��������: [1:0]���صȼ� 00:100% 01:50% 10:25% 11:12.5%  ���� 
 
    .o_recive_package       ( w_recive_package      )  , // �������ݰ��� 
    .o_recive_package_multi ( w_recive_package_multi)  , // �������ݰ�������
    .o_send_package         ( w_send_package        )  , // �������ݰ�����
    .o_send_package_multi   ( w_send_package_multi  )  , // �������ݰ���������
 
    .i_flow_data            ( w_flow_ctrl_input_data )  , // �˿����� (����ѡ���)
    .i_flow_data_keep       ( w_flow_ctrl_input_keep )  , // �˿����������ź� (����ѡ���)
    .i_flow_valid           ( w_flow_ctrl_input_valid)  , // �˿�������Ч (����ѡ���)
    .o_flow_ready           ( w_flow_ready           )  , // �˿����ݾ����ź�
    .i_flow_last            ( w_flow_ctrl_input_last )  , // ������������־ (����ѡ���)
 
    .o_flow_data            ( w_flow_data_out       )  , // ���غ�˿����� 
    .o_flow_data_keep       ( w_flow_data_keep_out  )  , // ���غ����������ź�
    .o_flow_valid           ( w_flow_valid_out      )  , // ���غ�������Ч
    .i_flow_ready           ( i_mac_axi_data_ready  )  , // ����ģ��ready�ź�
    .o_flow_last            ( w_flow_last_out       )    // ���غ����ݽ�����־

);

//-------------------- metadataƴ����� --------------------
always @(posedge i_clk) begin
    if (i_rst)
        ro_cross_metadata <= {METADATA_WIDTH{1'b0}};
    else
        ro_cross_metadata <= {
            ri_rtag_sequence      , // [80:65] R-TAG�ֶ� (16bit)
            ri_port_speed         , // [64:63] (2bit)
            ri_vlan_pri           , // [62:60] (3bit)
            ri_tx_prot            , // [59:52] tx_prot (8bit, �ں�ACLת���˿�)
            ri_acl_frmtype        , // [51:44] (8bit)
            ri_acl_cb_streamhandle, // [43:36] stream_handle (8bit)
            8'd0                  , // [35:28] �����ֶ� (8bit)
            ri_frm_vlan_flag      , // [27] (1bit)
            r_rx_port             , // [26:19] ����˿� (8bit)
            4'd0                  , // [18:15] ���� (4bit)
            ri_frm_cb_op          , // [14:13] [1]:rtag_flag [0]:cb_frm (2bit)
            w_discard             , // [12] ����λ (1bit)
            ri_frm_qbu            , // [11] (1bit)
            ri_timestamp_addr     , // [10:4] (7bit)
            4'd0                    // [3:0] ���� (4bit)

        };
end

//-------------------- metadata_valid�����߼� --------------------
// swlist_vld������־ 
always @(posedge i_clk) begin
    if (i_rst)
        r_swlist_vld_flag <= 1'b0;
    else
        r_swlist_vld_flag <= (w_both_vld_ready == 1'd1) ? 1'b0 : ((i_swlist_vld == 1'd1) ? 1'b1 : r_swlist_vld_flag);
end

// acl_vld������־  
always @(posedge i_clk) begin
    if (i_rst)
        r_acl_vld_flag <= 1'b0;
    else
        r_acl_vld_flag <= (w_both_vld_ready == 1'd1) ? 1'b0 : ((i_acl_vld == 1'd1) ? 1'b1 : r_acl_vld_flag);
end

// ����vld���Ѵ�����ָʾ�ź�
assign w_both_vld_ready = r_swlist_vld_flag == 1'd1 && r_acl_vld_flag == 1'd1 ? 1'd1 : 1'd0;

// metadata_valid��������ͬ���������ɺ�����������������
always @(posedge i_clk) begin
    if (i_rst)
        ro_cross_metadata_valid <= 1'b0;
    else
        ro_cross_metadata_valid <= (((w_flow_valid_out == 1'd1 && ro_mac_axi_data_valid == 1'd0) || (ro_mac_axi_data_valid == 1'd0 && r_fifo_rd_en == 1'd1 && r_need_flow_ctrl == 1'd0))) ? 1'd1  
                                   : 1'b0;
end

always @(posedge i_clk) begin
    if (i_rst)
        ro_cross_metadata_last <= 1'b0;
    else
        ro_cross_metadata_last <=  (((w_flow_valid_out == 1'd1 && ro_mac_axi_data_valid == 1'd0) || (ro_mac_axi_data_valid == 1'd0 && r_fifo_rd_en == 1'd1 && r_need_flow_ctrl == 1'd0))) ? 1'd1  
                                   : 1'b0;
end

always @(posedge i_clk) begin
    if (i_rst)
        ro_mac_port_axi_data <= {PORT_MNG_DATA_WIDTH{1'b0}};
    else
        ro_mac_port_axi_data <= (r_need_flow_ctrl == 1'd1) ? (w_flow_valid_out ? w_flow_data_out : {PORT_MNG_DATA_WIDTH{1'b0}}) :
                                (r_fifo_rd_en) ? w_fifo_out_data : {PORT_MNG_DATA_WIDTH{1'b0}};
end

always @(posedge i_clk) begin
    if (i_rst)
        ro_mac_axi_data_keep <= {(PORT_MNG_DATA_WIDTH/8){1'b0}};
    else
        ro_mac_axi_data_keep <= (r_need_flow_ctrl == 1'd1) ? (w_flow_valid_out ? w_flow_data_keep_out :{(PORT_MNG_DATA_WIDTH/8){1'b0}} ):
                                (r_fifo_rd_en == 1'd1) ? w_fifo_out_keep : {(PORT_MNG_DATA_WIDTH/8){1'b0}};
end

always @(posedge i_clk) begin
    if (i_rst)
        ro_mac_axi_data_valid <= 1'b0;
    else
        ro_mac_axi_data_valid <= (r_need_flow_ctrl == 1'd1) ? w_flow_valid_out : r_fifo_rd_en;
end

always @(posedge i_clk) begin
    if (i_rst)
        ro_mac_axi_data_last <= 1'b0;
    else
        ro_mac_axi_data_last <= (r_need_flow_ctrl == 1'd1) ? (w_flow_valid_out ? w_flow_last_out : 1'b0) :
                                (r_fifo_rd_en == 1'd1) ? w_fifo_out_last : 1'b0;
end

always @(posedge i_clk) begin
    if (i_rst)
        ro_mac_axi_data_user <= 16'd0;
    else
        ro_mac_axi_data_user <= r_frame_user;
end

// ���������
assign o_mac_port_axi_data          = ro_mac_port_axi_data                                     ;
assign o_mac_axi_data_keep          = ro_mac_axi_data_keep                                     ;
assign o_mac_axi_data_valid         = ro_mac_axi_data_valid                                    ;
assign o_mac_axi_data_last          = ro_mac_axi_data_last                                     ;
assign o_mac_axi_data_user          = ro_mac_axi_data_user                                     ;
assign o_mac_axi_data_ready         = ~w_fifo_full                                             ; // FIFOδ��ʱ���Խ�������

// metadata���
assign o_cross_metadata             = ro_cross_metadata                                        ;
assign o_cross_metadata_valid       = ro_cross_metadata_valid                                  ;
assign o_cross_metadata_last        = ro_cross_metadata_last                                   ;

// �������źţ���ʱ��Ĭ��ֵ����������չ��
assign o_port_rx_ultrashort_frm     = 1'b0                                                     ;
assign o_port_rx_overlength_frm     = 1'b0                                                     ;
// assign o_port_rx_crcerr_frm         = ri_mac_port_axi_data[CROSS_DATA_WIDTH]                   ; // ���λ��ʾCRC����
assign o_port_rx_loopback_frm_cnt   = 16'd0                                                    ;
assign o_port_broadflow_drop_cnt    = 16'd0                                                    ;
assign o_port_multiflow_drop_cnt    = 16'd0                                                    ;
assign o_port_diag_state            = {12'd0, w_send_package[3:0]}                             ; // ��4λ��ʾ���Ͱ�����
endmodule