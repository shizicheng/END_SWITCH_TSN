/*
 * ���ܣ�
 *  
 */

 
`timescale 1ns / 1ns
module rx_port_cache_mng#(
    parameter                                                           PORT_NUM                    = 8                         , // �������Ķ˿���
    parameter                                                           PORT_MNG_DATA_WIDTH         = 8                         , // Mac_port_mng ����λ��
    parameter                                                           METADATA_WIDTH              = 81                        , // ��Ϣ��λ��
    parameter                                                           CROSS_DATA_WIDTH            = 8                         , // �ۺ��������
    parameter                                                           PORT_FIFO_PRI_NUM           = 8                         , // ���ȼ�FIFO����
    parameter                                                           RAM_DEPTH                   = 1024                      , // RAM���
    parameter                                                           RAM_ADDR_WIDTH              = 10                        , // RAM��ַ���
    parameter                                                           FIFO_DEPTH                  = 512                      , // FIFO���
    parameter                                                           REQ_TIMEOUT_CNT             = 1250                      , // req��ʱ����ֵ(5us @ 250MHz)
    parameter                                                           TIMEOUT_CNT_WIDTH           = 11                         // ��ʱ������λ��
)(
    /*---------------------------------------- ʱ�Ӻ͸�λ -------------------------------------------*/
    input               wire                                            i_clk                               , // 250MHz
    input               wire                                            i_rst                               ,
    
    /*---------------------------------------- �����MAC������ -------------------------------------------*/
    input               wire   [PORT_MNG_DATA_WIDTH-1:0]                i_mac_axi_data                     , // �˿�������  
    input               wire   [(PORT_MNG_DATA_WIDTH/8)-1:0]            i_mac_axi_data_keep                , // �˿����������룬��Ч�ֽ�ָʾ
    input               wire                                            i_mac_axi_data_valid               , // �˿�������Ч
    output              wire                                            o_mac_axi_data_ready               , // �˿����ݾ����ź�,��ʾ��ǰģ��׼���ý�������
    input               wire                                            i_mac_axi_data_last                , // ������������ʶ
    input               wire   [15:0]                                   i_mac_axi_data_user                , // �Ƿ�ؼ�֡ + ���ĳ���
    
    /*---------------------------------------- �����metadata�� -------------------------------------------*/
    input               wire   [METADATA_WIDTH-1:0]                     i_cross_metadata                   , // ����metadata����
    input               wire                                            i_cross_metadata_valid             , // ����metadata������Ч�ź�
    input               wire                                            i_cross_metadata_last              , // ����metadata������ʶ
    output              wire                                            o_cross_metadata_ready             , // metadata��ѹ��ˮ��

    /*---------------------------------------- ������������ߵ������� -------------------------------------------*/ 

    output              wire   [15:0]                                   o_mac_cross_port_axi_user          , // �Ƿ�ؼ�֡ + ���ĳ���
    output              wire   [CROSS_DATA_WIDTH-1:0]                   o_mac_cross_port_axi_data          , // �˿������������λ��ʾcrcerr
    output              wire   [(CROSS_DATA_WIDTH/8)-1:0]               o_mac_cross_axi_data_keep          , // �˿����������룬��Ч�ֽ�ָʾ
    output              wire                                            o_mac_cross_axi_data_valid         , // �˿�������Ч
    input               wire                                            i_mac_cross_axi_data_ready         , // �������߾ۺϼܹ���ѹ��ˮ���ź�
    output              wire                                            o_mac_cross_axi_data_last          , // ������������ʶ
    
    /*---------------------------------------- ������������ߵ�metadata�� -------------------------------------------*/
    output              wire   [METADATA_WIDTH-1:0]                     o_cross_metadata                   , // �ۺ�����metadata����
    output              wire                                            o_cross_metadata_valid             , // �ۺ�����metadata������Ч�ź�
    output              wire                                            o_cross_metadata_last              , // ��Ϣ��������ʶ
    input               wire                                            i_cross_metadata_ready             , // ����ģ�鷴ѹ��ˮ��
    
    /*---------------------------------------- �� PORT �ؼ�֡��������� -------------------------------------------*/ 
    output              wire   [CROSS_DATA_WIDTH-1:0]                   o_emac_port_axi_data               , // �˿������������λ��ʾcrcerr
    output              wire   [15:0]                                   o_emac_port_axi_user               ,
    output              wire   [(CROSS_DATA_WIDTH/8)-1:0]               o_emac_axi_data_keep               , // �˿����������룬��Ч�ֽ�ָʾ
    output              wire                                            o_emac_axi_data_valid              , // �˿�������Ч
    input               wire                                            i_emac_axi_data_ready              , // �������߾ۺϼܹ���ѹ��ˮ���ź�
    output              wire                                            o_emac_axi_data_last               , // ������������ʶ
    /*---------------------------------------- �� PORT �ۺ���Ϣ�� -------------------------------------------*/
    output              wire   [METADATA_WIDTH-1:0]                     o_emac_metadata                    , // ���� metadata ����
    output              wire                                            o_emac_metadata_valid              , // ���� metadata ������Ч�ź�
    output              wire                                            o_emac_metadata_last               , // ��Ϣ��������ʶ
    input               wire                                            i_emac_metadata_ready              , // ����ģ�鷴ѹ��ˮ�� 
    
    /*---------------------------------------- �뷢�Ͷ˵�req-ack���� -------------------------------------------*/
    output              wire                                            o_rtag_flag                        , // �Ƿ�Я��rtag��ǩ,��CBҵ��֡,��Ҫ�ȹ�CBģ������Ƿ�����,������crossbar
    output              wire   [15:0]                                   o_rtag_squence                     , // rtag_squencenum
    output              wire   [7:0]                                    o_stream_handle                    , // ACL��ʶ��,��������ÿ��������ά���Լ���

    input               wire                                            i_pass_en                          , // �жϽ�������Խ��ո�֡
    input               wire                                            i_discard_en                       , // �жϽ�������Զ�����֡
    input               wire                                            i_judge_finish                     , // �жϽ������ʾ���α��ĵ��ж����

    output              wire                                            o_tx_req                           , // ���Ͷ˵�req�ź�
    input               wire                                            i_mac_tx0_ack                      , // �˿�0��Ӧʹ���ź�
    input               wire   [PORT_FIFO_PRI_NUM-1:0]                  i_mac_tx0_ack_rst                  , // �˿�0���ȼ��������
    input               wire                                            i_mac_tx1_ack                      , // �˿�1��Ӧʹ���ź�
    input               wire   [PORT_FIFO_PRI_NUM-1:0]                  i_mac_tx1_ack_rst                  , // �˿�1���ȼ��������  
    input               wire                                            i_mac_tx2_ack                      , // �˿�2��Ӧʹ���ź�
    input               wire   [PORT_FIFO_PRI_NUM-1:0]                  i_mac_tx2_ack_rst                  , // �˿�2���ȼ��������
    input               wire                                            i_mac_tx3_ack                      , // �˿�3��Ӧʹ���ź�
    input               wire   [PORT_FIFO_PRI_NUM-1:0]                  i_mac_tx3_ack_rst                  , // �˿�3���ȼ��������
    input               wire                                            i_mac_tx4_ack                      , // �˿�4��Ӧʹ���ź�
    input               wire   [PORT_FIFO_PRI_NUM-1:0]                  i_mac_tx4_ack_rst                  , // �˿�4���ȼ��������
    input               wire                                            i_mac_tx5_ack                      , // �˿�5��Ӧʹ���ź�
    input               wire   [PORT_FIFO_PRI_NUM-1:0]                  i_mac_tx5_ack_rst                  , // �˿�5���ȼ��������
    input               wire                                            i_mac_tx6_ack                      , // �˿�6��Ӧʹ���ź�
    input               wire   [PORT_FIFO_PRI_NUM-1:0]                  i_mac_tx6_ack_rst                  , // �˿�6���ȼ��������
    input               wire                                            i_mac_tx7_ack                      , // �˿�7��Ӧʹ���ź�
    input               wire   [PORT_FIFO_PRI_NUM-1:0]                  i_mac_tx7_ack_rst                  , // �˿�7���ȼ��������
    
    /*---------------------------------------- ƽ̨�Ĵ������� -------------------------------------------*/
    input               wire                                            i_port_rxmac_down_regs             , // �˿ڽ��շ���MAC�ر�ʹ��
    input               wire                                            i_port_broadcast_drop_regs         , // �˿ڹ㲥֡����ʹ��
    input               wire                                            i_port_multicast_drop_regs         , // �˿��鲥֡����ʹ��
    input               wire                                            i_port_loopback_drop_regs          , // �˿ڻ���֡����ʹ��
    input               wire   [47:0]                                   i_port_mac_regs                    , // �˿ڵ�MAC��ַ
    input               wire                                            i_port_mac_vld_regs                , // ʹ�ܶ˿�MAC��ַ��Ч
    input               wire   [15:0]                                   i_port_mtu_regs                    , // MTU����ֵ
    input               wire   [PORT_NUM-1:0]                           i_port_mirror_frwd_regs            , // ����ת���Ĵ���
    input               wire   [31:0]                                   i_port_flowctrl_cfg_regs           , // ������������
    input               wire   [15:0]                                   i_port_rx_ultrashortinterval_num   , // ֡���
    
    /*---------------------------------------- ACL�Ĵ��� -------------------------------------------*/
    input               wire   [2:0]                                    i_acl_port_sel                     , // ѡ��Ҫ���õĶ˿�
    input               wire                                            i_acl_clr_list_regs                , // ��ռĴ����б�
    output              wire                                            o_acl_list_rdy_regs                , // ���üĴ�����������
    input               wire   [9:0]                                    i_acl_item_sel_regs                , // ������Ŀѡ��
    input               wire   [5:0]                                    i_acl_item_waddr_regs              , // ÿ����Ŀ���֧�ֱȶ�64�ֽ�
    input               wire   [7:0]                                    i_acl_item_din_regs                , // ��Ҫ�Ƚϵ��ֽ�����
    input               wire                                            i_acl_item_we_regs                 , // ����ʹ���ź�
    input               wire   [15:0]                                   i_acl_item_rslt_regs               , // ƥ��Ľ��ֵ
    input               wire                                            i_acl_item_complete_regs           , // �˿�ACL�����������ʹ���ź�
    
    /*---------------------------------------- ״̬����ϼĴ��� -------------------------------------------*/
    output              wire   [31:0]                                   o_port_diag_state                  , // �˿�״̬�Ĵ���
    output              wire   [31:0]                                   o_port_rx_ultrashort_frm           , // �˿ڽ��ճ���֡
    output              wire   [31:0]                                   o_port_rx_overlength_frm           , // �˿ڽ��ճ���֡
    output              wire   [31:0]                                   o_port_rx_crcerr_frm               , // �˿ڽ���CRC����֡
    output              wire   [31:0]                                   o_port_rx_loopback_frm_cnt         , // �˿ڽ��ջ���֡������ֵ
    output              wire   [31:0]                                   o_port_broadflow_drop_cnt          , // �˿ڹ㲥��������֡������ֵ
    output              wire   [31:0]                                   o_port_multiflow_drop_cnt          , // �˿��鲥��������֡������ֵ
    output              wire   [63:0]                                   o_port_rx_byte_cnt                 , // �˿ڽ����ֽڸ���������ֵ
    output              wire   [31:0]                                   o_port_rx_frame_cnt                  // �˿ڽ���֡����������ֵ
);

/*---------------------------------------- �ڲ��������� -------------------------------------------*/
localparam                  QUEUE_SIZE              = 32                                                    ; // �����������
localparam                  QUEUE_ADDR_WIDTH        = 5                                                     ; // ���е�ַλ��
localparam                  FRAME_INFO_WIDTH        = METADATA_WIDTH + 16                                   ; // ֡��Ϣλ��(metadata + user)
localparam                  TIMEOUT_CNT_MAX         = REQ_TIMEOUT_CNT - 1                                   ; // ��ʱ�������ֵ

/*---------------------------------------- �ڲ��Ĵ������������� -------------------------------------------*/

// ��������ź�
reg                                     ri_mac_axi_data_valid          ;
reg    [PORT_MNG_DATA_WIDTH-1:0]        ri_mac_axi_data                ;
reg    [(PORT_MNG_DATA_WIDTH/8)-1:0]    ri_mac_axi_data_keep           ;
reg                                     ri_mac_axi_data_last           ;
reg    [15:0]                           ri_mac_axi_data_user           ;
reg                                     ri_cross_metadata_valid        ; 
reg                                     ri_cross_metadata_valid_1d     ;
reg    [METADATA_WIDTH-1:0]             ri_cross_metadata              ;
reg                                     ri_cross_metadata_last         ;
reg                                     ri_pass_en                     ;
reg                                     ri_discard_en                  ;
reg                                     ri_judge_finish                ;
reg                                     ri_mac_tx0_ack                 ;
reg    [PORT_FIFO_PRI_NUM-1:0]          ri_mac_tx0_ack_rst             ;
reg                                     ri_mac_tx1_ack                 ;
reg    [PORT_FIFO_PRI_NUM-1:0]          ri_mac_tx1_ack_rst             ;
reg                                     ri_mac_tx2_ack                 ;
reg    [PORT_FIFO_PRI_NUM-1:0]          ri_mac_tx2_ack_rst             ;
reg                                     ri_mac_tx3_ack                 ;
reg    [PORT_FIFO_PRI_NUM-1:0]          ri_mac_tx3_ack_rst             ;
reg                                     ri_mac_tx4_ack                 ;
reg    [PORT_FIFO_PRI_NUM-1:0]          ri_mac_tx4_ack_rst             ;
reg                                     ri_mac_tx5_ack                 ;
reg    [PORT_FIFO_PRI_NUM-1:0]          ri_mac_tx5_ack_rst             ;
reg                                     ri_mac_tx6_ack                 ;
reg    [PORT_FIFO_PRI_NUM-1:0]          ri_mac_tx6_ack_rst             ;
reg                                     ri_mac_tx7_ack                 ;
reg    [PORT_FIFO_PRI_NUM-1:0]          ri_mac_tx7_ack_rst             ;

// ����Ĵ���
reg                                     ro_mac_axi_data_ready          ;
reg                                     ro_cross_metadata_ready        ;
reg    [15:0]                           ro_mac_cross_port_axi_user     ;
reg    [CROSS_DATA_WIDTH-1:0]           ro_mac_cross_port_axi_data     ;
reg    [(CROSS_DATA_WIDTH/8)-1:0]       ro_mac_cross_axi_data_keep     ;
reg                                     ro_mac_cross_axi_data_valid    ;
reg                                     ro_mac_cross_axi_data_valid_d1 ;
reg                                     ro_mac_cross_axi_data_last     ;
reg    [METADATA_WIDTH-1:0]             ro_cross_metadata              ;
reg                                     ro_cross_metadata_valid        ;
reg                                     ro_cross_metadata_last         ;
reg                                     ro_rtag_flag                   ;
reg    [15:0]                           ro_rtag_squence                ;
reg    [7:0]                            ro_stream_handle               ;
reg                                     ro_tx_req                      ;
reg                                     ro_tx_req_d1                   ;

// ���й�����ؼĴ���
reg    [QUEUE_ADDR_WIDTH-1:0]           r_wr_addr                      ; // д��ַ
reg    [QUEUE_ADDR_WIDTH-1:0]           r_rd_addr                      ; // ����ַ
reg    [QUEUE_ADDR_WIDTH:0]             r_ram_data_cnt                 ; // FIFO����
reg                                     r_queue_full                   ; // ��������־
reg                                     r_queue_empty                  ; // ���пձ�־

// ����RAM����ź�
wire   [RAM_ADDR_WIDTH-1:0]             w_data_ram_wr_addr             ;
wire   [RAM_ADDR_WIDTH-1:0]             w_data_ram_rd_addr             ;
wire   [PORT_MNG_DATA_WIDTH + (PORT_MNG_DATA_WIDTH/8)-1:0] w_data_ram_wr_data ;
wire   [PORT_MNG_DATA_WIDTH + (PORT_MNG_DATA_WIDTH/8)-1:0] w_data_ram_rd_data ;
wire                                    w_data_ram_we                  ;
wire                                    w_data_ram_re                  ;

// ��ϢRAM����ź�
wire   [QUEUE_ADDR_WIDTH-1:0]           w_info_ram_wr_addr             ;
wire   [QUEUE_ADDR_WIDTH-1:0]           w_info_ram_rd_addr             ;
wire   [FRAME_INFO_WIDTH-1:0]           w_info_ram_wr_data             ;
wire   [FRAME_INFO_WIDTH-1:0]           w_info_ram_rd_data             ;
wire                                    w_info_ram_we                  ;
reg                                     r_info_ram_we                  ; 
reg                                     r_info_ram_re                  ;

// ֡������ؼĴ���
wire                                    w_frame_read_end               ;
reg                                     r_frame_writing                ; // ֡д���־
reg                                     r_frame_reading                ; // ֡��ȡ��־
reg    [RAM_ADDR_WIDTH-1:0]             r_current_frame_start_addr     ; // ��ǰ֡��ʼ��ַ
reg    [RAM_ADDR_WIDTH-1:0]             r_current_frame_end_addr       ; // ��ǰ֡������ַ
reg    [RAM_ADDR_WIDTH-1:0]             r_frame_start_addrs [QUEUE_SIZE-1:0] ; // ÿ���������Ӧ��֡��ʼ��ַ
reg    [RAM_ADDR_WIDTH-1:0]             r_frame_end_addrs   [QUEUE_SIZE-1:0] ; // ÿ���������Ӧ��֡������ַ
reg    [RAM_ADDR_WIDTH-1:0]             r_data_wr_ptr                  ; // ����RAMдָ��
reg    [RAM_ADDR_WIDTH-1:0]             r_data_ram_rd_ptr              ; // ����RAM��ָ��

// metadata������ؼĴ���
reg                                     r_rtag_flag                    ; // rtag��־λ
reg    [15:0]                           r_rtag_squence                 ; // rtag���к�
reg    [7:0]                            r_stream_handle                ; // �����
reg    [2:0]                            r_vlan_pri                     ; // VLAN���ȼ�

// ��ǰ����֡�Ƿ�Ϊ�ؼ�֡
reg                                     r_current_is_critical          ;

// CB������ؼĴ���
reg                                     r_cb_processing                ; // CB�����б�־
reg                                     r_cb_req_sent                  ; // CB�����ѷ��ͱ�־
reg                                     r_cb_result_rcvd               ; // CB����ѽ��ձ�־
reg                                     r_pass_result                  ; // ͨ�����

// req-ack������ؼĴ���
reg                                     r_req_sent                     ; // req�ѷ��ͱ�־
reg    [TIMEOUT_CNT_WIDTH-1:0]          r_timeout_cnt                  ; // ��ʱ������
reg                                     r_timeout_flag                 ; // ��ʱ��־
reg    [PORT_NUM-1:0]                   r_ack_received                 ; // ACK���ձ�־
reg    [PORT_NUM-1:0]                   r_ack_expected                 ; // ������ACK

// ���ȼ�������ؼĴ���
reg    [QUEUE_ADDR_WIDTH-1:0]           r_current_process_addr         ; // ��ǰ�����ַ
reg                                     r_process_complete             ; // ������ɱ�־
reg    [2:0]                            r_frame_pri         [QUEUE_SIZE-1:0] ; // ÿ������������ȼ���3λVLAN���ȼ���
reg                                     r_frame_valid       [QUEUE_SIZE-1:0] ; // ÿ�����������Ч��־
reg                                     r_frame_end_addr_valid [QUEUE_SIZE-1:0] ; // ÿ��������Ľ�����ַ��Ч��־
// two-stage register for r_info_ram_re
reg                                     r_info_ram_re_d1               ;
reg                                     r_info_ram_re_d2               ;
reg                                     r_process_complete_d1          ;
// ���ȼ�ѡ���ź�
wire   [2:0]                            r_max_pri                      ; // ������ȼ�ֵ
wire   [QUEUE_ADDR_WIDTH-1:0]           r_next_addr                    ; // ��һ�������ַ

wire                                    w_tx_req                       ;
wire                                    w_recivedall_ack               ;

reg    [15:0]                           r_data_out_cnt                 ;
reg    [15:0]                           r_data_out_len                 ;

wire   [METADATA_WIDTH-1:0]             w_current_metadata             ;
// ״̬��־
// reg                         r_input_ready                                                          ; // ���������־
// reg                         r_output_valid                                                         ; // �����Ч��־


assign w_recivedall_ack = ((r_ack_received & r_ack_expected) == r_ack_expected) && (r_ack_expected != {PORT_NUM{1'b0}}) ? 1'd1 : 1'd0;

assign w_frame_read_end = (o_mac_cross_axi_data_valid == 1'b1) && (o_mac_cross_axi_data_last == 1'b1) ? 1'd1 : 1'd0 ;

// �ؼ�֡�жϣ�user�ź����λ��metadata[11]
wire   w_is_critical_frame;
assign w_is_critical_frame = (((w_current_metadata[11] == 1'b1) || (w_info_ram_rd_data[15] == 1'b1)) && (w_current_metadata[13] == 1'b1))? 1'd1 : 1'd0 ;

 

/*---------------------------------------- �����źŴ��� -------------------------------------------*/
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        ri_mac_axi_data_valid      <= 1'b0;
        ri_mac_axi_data            <= {PORT_MNG_DATA_WIDTH{1'b0}};
        ri_mac_axi_data_keep       <= {(PORT_MNG_DATA_WIDTH/8){1'b0}};
        ri_mac_axi_data_last       <= 1'b0;
        ri_mac_axi_data_user       <= 16'b0;
        ri_cross_metadata_valid    <= 1'b0;
        ri_cross_metadata_valid_1d <= 1'b0;
        ri_cross_metadata          <= {METADATA_WIDTH{1'b0}};
        ri_cross_metadata_last     <= 1'b0;
        ri_pass_en                 <= 1'b0;
        ri_discard_en              <= 1'b0;
        ri_judge_finish            <= 1'b0;
        ri_mac_tx0_ack             <= 1'b0;
        ri_mac_tx0_ack_rst         <= {PORT_FIFO_PRI_NUM{1'b0}};
        ri_mac_tx1_ack             <= 1'b0;
        ri_mac_tx1_ack_rst         <= {PORT_FIFO_PRI_NUM{1'b0}};
        ri_mac_tx2_ack             <= 1'b0;
        ri_mac_tx2_ack_rst         <= {PORT_FIFO_PRI_NUM{1'b0}};
        ri_mac_tx3_ack             <= 1'b0;
        ri_mac_tx3_ack_rst         <= {PORT_FIFO_PRI_NUM{1'b0}};
        ri_mac_tx4_ack             <= 1'b0;
        ri_mac_tx4_ack_rst         <= {PORT_FIFO_PRI_NUM{1'b0}};
        ri_mac_tx5_ack             <= 1'b0;
        ri_mac_tx5_ack_rst         <= {PORT_FIFO_PRI_NUM{1'b0}};
        ri_mac_tx6_ack             <= 1'b0;
        ri_mac_tx6_ack_rst         <= {PORT_FIFO_PRI_NUM{1'b0}};
        ri_mac_tx7_ack             <= 1'b0;
        ri_mac_tx7_ack_rst         <= {PORT_FIFO_PRI_NUM{1'b0}};
    end else begin
        ri_mac_axi_data_valid      <= i_mac_axi_data_valid;
        ri_mac_axi_data            <= i_mac_axi_data;
        ri_mac_axi_data_keep       <= i_mac_axi_data_keep;
        ri_mac_axi_data_last       <= i_mac_axi_data_last;
        ri_mac_axi_data_user       <= i_mac_axi_data_user;
        ri_cross_metadata_valid    <= i_cross_metadata_valid;
        ri_cross_metadata_valid_1d <= ri_cross_metadata_valid;
        ri_cross_metadata          <= i_cross_metadata;
        ri_cross_metadata_last     <= i_cross_metadata_last;
        ri_pass_en                 <= i_pass_en;
        ri_discard_en              <= i_discard_en;
        ri_judge_finish            <= i_judge_finish;
        ri_mac_tx0_ack             <= i_mac_tx0_ack;
        ri_mac_tx0_ack_rst         <= i_mac_tx0_ack_rst;
        ri_mac_tx1_ack             <= i_mac_tx1_ack;
        ri_mac_tx1_ack_rst         <= i_mac_tx1_ack_rst;
        ri_mac_tx2_ack             <= i_mac_tx2_ack;
        ri_mac_tx2_ack_rst         <= i_mac_tx2_ack_rst;
        ri_mac_tx3_ack             <= i_mac_tx3_ack;
        ri_mac_tx3_ack_rst         <= i_mac_tx3_ack_rst;
        ri_mac_tx4_ack             <= i_mac_tx4_ack;
        ri_mac_tx4_ack_rst         <= i_mac_tx4_ack_rst;
        ri_mac_tx5_ack             <= i_mac_tx5_ack;
        ri_mac_tx5_ack_rst         <= i_mac_tx5_ack_rst;
        ri_mac_tx6_ack             <= i_mac_tx6_ack;
        ri_mac_tx6_ack_rst         <= i_mac_tx6_ack_rst;
        ri_mac_tx7_ack             <= i_mac_tx7_ack;
        ri_mac_tx7_ack_rst         <= i_mac_tx7_ack_rst;
    end
end

/*---------------------------------------- ���й����߼� -------------------------------------------*/
// ������֡������
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_ram_data_cnt <= {(QUEUE_ADDR_WIDTH+1){1'b0}};
    end else begin
        r_ram_data_cnt <= ((ri_cross_metadata_valid == 1'b1) && (r_queue_full == 1'b0) && !((r_process_complete == 1'b1) && (r_queue_empty == 1'b0))) ? 
                        (r_ram_data_cnt + {{QUEUE_ADDR_WIDTH{1'b0}}, 1'b1}) :
                      ((r_process_complete == 1'b1) && (r_queue_empty == 1'b0) && !((ri_cross_metadata_valid == 1'b1) && (r_queue_full == 1'b0))) ? 
                        (r_ram_data_cnt - {{QUEUE_ADDR_WIDTH{1'b0}}, 1'b1}) :
                      r_ram_data_cnt;
    end
end

// ������/�ձ�־
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_queue_full <= 1'b0;
    end else begin
        r_queue_full <= (r_ram_data_cnt[QUEUE_ADDR_WIDTH] == 1'b1) ? 1'b1 : 1'b0;
    end
end

always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_queue_empty <= 1'b1;
    end else begin
        r_queue_empty <= (r_ram_data_cnt == {(QUEUE_ADDR_WIDTH+1){1'b0}}) ? 1'b1 : 1'b0;
    end
end

// д��ַ����
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_wr_addr <= {QUEUE_ADDR_WIDTH{1'b0}};
    end else begin
        r_wr_addr <= ri_mac_axi_data_last == 1'd1 && ri_mac_axi_data_valid == 1'b1 && r_queue_full == 1'b0 && (r_wr_addr == (QUEUE_SIZE - {{(QUEUE_ADDR_WIDTH-1){1'b0}},1'b1})) ? {QUEUE_ADDR_WIDTH{1'b0}} : 
                     ri_mac_axi_data_last == 1'd1 && ri_mac_axi_data_valid == 1'b1 && r_queue_full == 1'b0 ? (r_wr_addr + {{(QUEUE_ADDR_WIDTH-1){1'b0}}, 1'b1}) :
                     r_wr_addr;
    end
end

// ����ַ���� - �������ȼ�ѡ��������
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_rd_addr <= {QUEUE_ADDR_WIDTH{1'b0}};
    end else begin
        r_rd_addr <= r_info_ram_we == 1'b1 ? r_next_addr : r_rd_addr;
    end
end

/*---------------------------------------- ����RAMд����� -------------------------------------------*/
// ����RAMдָ��
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_data_wr_ptr <= {RAM_ADDR_WIDTH{1'b0}};
    end else begin
        r_data_wr_ptr <= ((ri_mac_axi_data_valid == 1'b1) && (ro_mac_axi_data_ready == 1'b1)) ?
                         ((r_data_wr_ptr == (RAM_DEPTH - 1)) ? {RAM_ADDR_WIDTH{1'b0}} : (r_data_wr_ptr + {{(RAM_ADDR_WIDTH-1){1'b0}}, 1'b1})) :
                         r_data_wr_ptr;
    end
end

// ֡д���־
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_frame_writing <= 1'b0;
    end else begin
        r_frame_writing <= ((ri_mac_axi_data_valid == 1'b1) && (ro_mac_axi_data_ready == 1'b1) && (r_frame_writing == 1'b0)) ? 1'b1 :
                          (((ri_mac_axi_data_valid == 1'b1) && (ri_mac_axi_data_last == 1'b1) && (ro_mac_axi_data_ready == 1'b1)) ? 1'b0 : r_frame_writing);
    end
end

// ��ǰ֡��ʼ��ַ
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_current_frame_start_addr <= {RAM_ADDR_WIDTH{1'b0}};
    end else begin
        r_current_frame_start_addr <= ((ri_mac_axi_data_valid == 1'b1) && (ro_mac_axi_data_ready == 1'b1) && (r_frame_writing == 1'b0)) ?
                                      r_data_wr_ptr : r_current_frame_start_addr;
    end
end

// ��ǰ֡������ַ
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_current_frame_end_addr <= {RAM_ADDR_WIDTH{1'b0}};
    end else begin
        r_current_frame_end_addr <= ((i_mac_axi_data_valid == 1'b1) && (i_mac_axi_data_last == 1'b1) && (ro_mac_axi_data_ready == 1'b1)) ?
                                    r_data_wr_ptr + 1'd1 : r_current_frame_end_addr;
    end
end

// �洢ÿ���������֡��ַ��Ϣ�����ȼ�����Ч��־
genvar gi;
generate
    for (gi = 0; gi < QUEUE_SIZE; gi = gi + 1) begin: g_queue_item
        always @(posedge i_clk) begin
            if (i_rst == 1'b1) begin
                r_frame_valid[gi]           <= 1'b0;
                r_frame_pri[gi]             <= 3'b0;
                r_frame_start_addrs[gi]     <= {RAM_ADDR_WIDTH{1'b0}};
            end else begin
                // ��д��֡ʱ����¼��ַ�����ȼ���������Ч��־
                r_frame_start_addrs[gi]     <= ((ri_cross_metadata_valid == 1'b1) && (r_queue_full == 1'b0) && (r_wr_addr == gi[QUEUE_ADDR_WIDTH-1:0])) ? r_data_wr_ptr : r_frame_start_addrs[gi];
                r_frame_pri[gi]             <= ((ri_cross_metadata_valid == 1'b1) && (r_queue_full == 1'b0) && (r_wr_addr == gi[QUEUE_ADDR_WIDTH-1:0])) ? ri_cross_metadata[62:60] : r_frame_pri[gi]; // VLAN���ȼ�λ
                r_frame_valid[gi]           <= ((r_process_complete == 1'b1) && (r_queue_empty == 1'b0) && (r_current_process_addr == gi[QUEUE_ADDR_WIDTH-1:0])) ? 1'b0 :
                                               ((ri_cross_metadata_valid == 1'b1) && (r_queue_full == 1'b0) && (r_wr_addr == gi[QUEUE_ADDR_WIDTH-1:0])) ? 1'b1 :  r_frame_valid[gi];
            end
        end
        
        // ��������֡������ַ����Ч��־
        always @(posedge i_clk) begin
            if (i_rst == 1'b1) begin
                r_frame_end_addrs[gi]       <= {RAM_ADDR_WIDTH{1'b0}};
                r_frame_end_addr_valid[gi]  <= 1'b0;
            end else begin
                // ֡���ݽ������ʱ����¼������ַ��������Ч��־
                r_frame_end_addrs[gi]       <= ((ri_mac_axi_data_valid == 1'd1) && (ri_mac_axi_data_last == 1'd1) && (r_queue_full == 1'b0) && (r_wr_addr == gi[QUEUE_ADDR_WIDTH-1:0])) ? r_current_frame_end_addr : r_frame_end_addrs[gi];
                r_frame_end_addr_valid[gi]  <= ((ri_mac_axi_data_valid == 1'd1) && (ri_mac_axi_data_last == 1'd1) && (r_queue_full == 1'b0) && (r_wr_addr == gi[QUEUE_ADDR_WIDTH-1:0])) ? 1'b1 :
                                               ((r_process_complete == 1'b1) && (r_queue_empty == 1'b0) && (r_current_process_addr == gi[QUEUE_ADDR_WIDTH-1:0])) ? 1'b0 : r_frame_end_addr_valid[gi];
            end
        end
    end
endgenerate

/*---------------------------------------- metadata���� -------------------------------------------*/
// ����metadata��RAM�е�λ�� (metadataλ�ڸ�λ��userλ�ڵ�15λ)
assign w_current_metadata = w_info_ram_rd_data[FRAME_INFO_WIDTH-1:16];

// rtag��־���� - �ӵ�ǰ���ж�ȡ��metadata����
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_rtag_flag <= 1'b0;
    end else begin
        r_rtag_flag <= (r_info_ram_re_d1 == 1'd1) ? w_current_metadata[14] : (r_process_complete == 1'b1) ? 1'b0 :r_rtag_flag;
    end
end

// ��ǰ����֡�Ƿ�Ϊ�ؼ�֡
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_current_is_critical <= 1'b0;
    end else begin
        r_current_is_critical <=  (r_process_complete == 1'b1) ? 1'b0 :
                                  (r_info_ram_re_d1 == 1'd1) ? w_is_critical_frame : 
                                  r_current_is_critical;
    end
end

// rtag���кŽ��� - �ӵ�ǰ���ж�ȡ��metadata����
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_rtag_squence <= 16'b0;
    end else begin
        r_rtag_squence <= (r_info_ram_re_d1 == 1'd1) ? w_current_metadata[80:65] : (r_process_complete == 1'b1) ? 1'b0 :r_rtag_squence;
    end
end

// ��������� - �ӵ�ǰ���ж�ȡ��metadata����
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_stream_handle <= 8'b0;
    end else begin
        r_stream_handle <= (r_info_ram_re_d1 == 1'd1) ? w_current_metadata[43:36] : (r_process_complete == 1'b1) ? 1'b0 :r_stream_handle;
    end
end

// VLAN���ȼ����� - �ӵ�ǰ���ж�ȡ��metadata����  
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_vlan_pri <= 3'b0;
    end else begin
        r_vlan_pri <= (r_info_ram_re_d1 == 1'd1) ? w_current_metadata[62:60] : (r_process_complete == 1'b1) ? 1'b0 :r_vlan_pri;
    end
end

/*---------------------------------------- CB�����߼� -------------------------------------------*/
// CB�����б�־
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_cb_processing <= 1'b0;
    end else begin
        r_cb_processing <= (r_rtag_flag == 1'b1 && r_queue_empty == 1'b0 && r_cb_processing == 1'd0 && r_cb_result_rcvd == 1'd0) ? 1'b1 :
                          ((ri_judge_finish == 1'b1) ? 1'b0 : r_cb_processing);
    end
end

// CB�����ѷ��ͱ�־
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_cb_req_sent <= 1'b0;
    end else begin
        r_cb_req_sent <= (r_cb_processing == 1'b1 && r_cb_req_sent == 1'b0 && r_cb_result_rcvd == 1'd0) ? 1'b1 : (ri_judge_finish == 1'b1) ? 1'b0 : r_cb_req_sent;
    end
end

// CB����ѽ��ձ�־
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_cb_result_rcvd <= 1'b0;
    end else begin
        r_cb_result_rcvd <= (r_cb_req_sent == 1'd1 && r_cb_result_rcvd == 1'b0) ? 1'b1 :
                           ((r_process_complete == 1'b1) ? 1'b0 : r_cb_result_rcvd);
    end
end

// ͨ�����
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_pass_result <= 1'b0;
    end else begin
        r_pass_result <= ((ri_judge_finish == 1'b1) && (ri_pass_en == 1'b1)) ? 1'b1 :
                        (((ri_judge_finish == 1'b1) && (ri_discard_en == 1'b1)) || r_process_complete == 1'd1 ? 1'b0 : r_pass_result);
    end
end

/*---------------------------------------- req-ack�����߼� -------------------------------------------*/
// req�ѷ��ͱ�־
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_req_sent <= 1'b0;
    end else begin
        r_req_sent <= (r_current_is_critical == 1'b0) && (ro_mac_cross_axi_data_valid_d1== 1'b1 || r_timeout_flag == 1'd1) ? 1'b0 :
                      ((r_current_is_critical == 1'b0) && (((r_info_ram_re_d2 == 1'd1) && (r_rtag_flag == 1'b0) && (r_queue_empty == 1'b0) && (r_req_sent == 1'b0)) ||
                      ((r_rtag_flag == 1'b1) && (r_cb_result_rcvd == 1'b1) && (r_pass_result == 1'b1) && (r_req_sent == 1'b0))))  ? 1'b1 :
                      r_req_sent;
    end
end

// ��ʱ������
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_timeout_cnt <= {TIMEOUT_CNT_WIDTH{1'b0}};
    end else begin
        r_timeout_cnt <=   (r_current_is_critical == 1'b0) && r_frame_reading == 1'd0 && r_req_sent == 1'b1  ?
                         ((r_timeout_cnt == TIMEOUT_CNT_MAX ) ? {TIMEOUT_CNT_WIDTH{1'b0}} : (r_timeout_cnt + {{(TIMEOUT_CNT_WIDTH-1){1'b0}}, 1'b1})) :
                         ((w_recivedall_ack == 1'b1) ? {TIMEOUT_CNT_WIDTH{1'b0}} : {TIMEOUT_CNT_WIDTH{1'b0}});
    end
end

// ��ʱ��־
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_timeout_flag <= 1'b0;
    end else begin
        r_timeout_flag <= (r_timeout_cnt == TIMEOUT_CNT_MAX) ? 1'b1 :  1'b0;
    end
end

/*---------------------------------------- ��������ź� -------------------------------------------*/
// ����������ؼ�֡��·ʱ������emac��ѹ���ƣ������ɶ����Ƿ�������
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        ro_mac_axi_data_ready <= 1'b0;
    end else begin
        ro_mac_axi_data_ready <= (r_queue_full == 1'b0) ? 1'b1 : 1'b0;
    end
end

// metadata�������ؼ�֡��·ʱ������emac��ѹ���ƣ������ɶ����Ƿ�������
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        ro_cross_metadata_ready <= 1'b0;
    end else begin
        ro_cross_metadata_ready <= (r_queue_full == 1'b0) ? 1'b1 : 1'b0;
    end
end

/*---------------------------------------- CB����ź� -------------------------------------------*/
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        ro_rtag_flag <= 1'b0;
    end else begin
        ro_rtag_flag <= ((r_cb_processing == 1'b1) && (r_cb_req_sent == 1'b0)) ? 1'b1 : 1'b0;
    end
end

always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        ro_rtag_squence <= 16'b0;
    end else begin
        ro_rtag_squence <= ((r_cb_processing == 1'b1) && (r_cb_req_sent == 1'b0)) ? 
                           w_current_metadata[80:65] : 16'b0;
    end
end

always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        ro_stream_handle <= 8'b0;
    end else begin
        ro_stream_handle <= ((r_cb_processing == 1'b1) && (r_cb_req_sent == 1'b0)) ? 
                            w_current_metadata[43:36] : 8'b0;
    end
end

/*---------------------------------------- ���ȼ�ѡ���߼� -------------------------------------------*/
// ���ȼ�ѡ������߼���ʹ�ö������ȽϽṹ��ѡ�����ȼ���ߵ���Ч������
// ���ж��ͬ���ȼ�֡��ѡ��������ӵģ�������С�ģ�

// ��һ���Ƚϣ������Ƚϣ�
wire   [2:0]                pri_cmp_l1      [15:0]                                              ; // ��һ�����ȼ��ȽϽ��
wire   [QUEUE_ADDR_WIDTH-1:0]           addr_cmp_l1     [15:0]                                  ; // ��һ����ַ�ȽϽ��
wire                        valid_cmp_l1    [15:0]                                              ; // ��һ����Ч��־�ȽϽ��

genvar gj;
generate
    for (gj = 0; gj < 16; gj = gj + 1) begin: g_pri_cmp_l1
        assign valid_cmp_l1[gj] = r_frame_valid[gj*2] | r_frame_valid[gj*2+1];
        assign pri_cmp_l1[gj]   = (!r_frame_valid[gj*2] && r_frame_valid[gj*2+1]) ? r_frame_pri[gj*2+1] :
                                  (r_frame_valid[gj*2] && !r_frame_valid[gj*2+1]) ? r_frame_pri[gj*2] :
                                  (r_frame_valid[gj*2] && r_frame_valid[gj*2+1]) ? 
                                  ((r_frame_pri[gj*2] > r_frame_pri[gj*2+1]) ? r_frame_pri[gj*2] : r_frame_pri[gj*2+1]) :
                                  3'b000;
        assign addr_cmp_l1[gj]  = (!r_frame_valid[gj*2] && r_frame_valid[gj*2+1]) ? (gj*2+1) :
                                  (r_frame_valid[gj*2] && !r_frame_valid[gj*2+1]) ? (gj*2) :
                                  (r_frame_valid[gj*2] && r_frame_valid[gj*2+1]) ? 
                                  ((r_frame_pri[gj*2] > r_frame_pri[gj*2+1]) ? (gj*2) : 
                                   (r_frame_pri[gj*2] < r_frame_pri[gj*2+1]) ? (gj*2+1) : (gj*2)) :
                                  {QUEUE_ADDR_WIDTH{1'b0}};
    end
endgenerate

// �ڶ����Ƚϣ�8���Ƚ�����
wire   [2:0]                pri_cmp_l2      [7:0]                                                          ; // �ڶ������ȼ��ȽϽ��
wire   [QUEUE_ADDR_WIDTH-1:0]           addr_cmp_l2     [7:0]                                   ; // �ڶ�����ַ�ȽϽ��
wire                        valid_cmp_l2    [7:0]                                                          ; // �ڶ�����Ч��־�ȽϽ��

generate
    for (gj = 0; gj < 8; gj = gj + 1) begin: g_pri_cmp_l2
        assign valid_cmp_l2[gj] = valid_cmp_l1[gj*2] | valid_cmp_l1[gj*2+1];
        assign pri_cmp_l2[gj]   = (!valid_cmp_l1[gj*2] && valid_cmp_l1[gj*2+1]) ? pri_cmp_l1[gj*2+1] :
                                  (valid_cmp_l1[gj*2] && !valid_cmp_l1[gj*2+1]) ? pri_cmp_l1[gj*2] :
                                  (valid_cmp_l1[gj*2] && valid_cmp_l1[gj*2+1]) ? 
                                  ((pri_cmp_l1[gj*2] > pri_cmp_l1[gj*2+1]) ? pri_cmp_l1[gj*2] : pri_cmp_l1[gj*2+1]) :
                                  3'b000;
        assign addr_cmp_l2[gj]  = (!valid_cmp_l1[gj*2] && valid_cmp_l1[gj*2+1]) ? addr_cmp_l1[gj*2+1] :
                                  (valid_cmp_l1[gj*2] && !valid_cmp_l1[gj*2+1]) ? addr_cmp_l1[gj*2] :
                                  (valid_cmp_l1[gj*2] && valid_cmp_l1[gj*2+1]) ? 
                                  ((pri_cmp_l1[gj*2] > pri_cmp_l1[gj*2+1]) ? addr_cmp_l1[gj*2] : 
                                   (pri_cmp_l1[gj*2] < pri_cmp_l1[gj*2+1]) ? addr_cmp_l1[gj*2+1] : addr_cmp_l1[gj*2]) :
                                  {QUEUE_ADDR_WIDTH{1'b0}};
    end
endgenerate

// �������Ƚϣ�4���Ƚ�����
wire   [2:0]                pri_cmp_l3      [3:0]                                                          ; // ���������ȼ��ȽϽ��
wire   [QUEUE_ADDR_WIDTH-1:0]           addr_cmp_l3     [3:0]                                   ; // ��������ַ�ȽϽ��
wire                        valid_cmp_l3    [3:0]                                                          ; // ��������Ч��־�ȽϽ��

generate
    for (gj = 0; gj < 4; gj = gj + 1) begin: g_pri_cmp_l3
        assign valid_cmp_l3[gj] = valid_cmp_l2[gj*2] | valid_cmp_l2[gj*2+1];
        assign pri_cmp_l3[gj]   = (!valid_cmp_l2[gj*2] && valid_cmp_l2[gj*2+1]) ? pri_cmp_l2[gj*2+1] :
                                  (valid_cmp_l2[gj*2] && !valid_cmp_l2[gj*2+1]) ? pri_cmp_l2[gj*2] :
                                  (valid_cmp_l2[gj*2] && valid_cmp_l2[gj*2+1]) ? 
                                  ((pri_cmp_l2[gj*2] > pri_cmp_l2[gj*2+1]) ? pri_cmp_l2[gj*2] : pri_cmp_l2[gj*2+1]) :
                                  3'b000;
        assign addr_cmp_l3[gj]  = (!valid_cmp_l2[gj*2] && valid_cmp_l2[gj*2+1]) ? addr_cmp_l2[gj*2+1] :
                                  (valid_cmp_l2[gj*2] && !valid_cmp_l2[gj*2+1]) ? addr_cmp_l2[gj*2] :
                                  (valid_cmp_l2[gj*2] && valid_cmp_l2[gj*2+1]) ? 
                                  ((pri_cmp_l2[gj*2] > pri_cmp_l2[gj*2+1]) ? addr_cmp_l2[gj*2] : 
                                   (pri_cmp_l2[gj*2] < pri_cmp_l2[gj*2+1]) ? addr_cmp_l2[gj*2+1] : addr_cmp_l2[gj*2]) :
                                  {QUEUE_ADDR_WIDTH{1'b0}};
    end
endgenerate

// ���ļ��Ƚϣ�2���Ƚ�����
wire   [2:0]                pri_cmp_l4      [1:0]                                                          ; // ���ļ����ȼ��ȽϽ��
wire   [QUEUE_ADDR_WIDTH-1:0]           addr_cmp_l4     [1:0]                                   ; // ���ļ���ַ�ȽϽ��
wire                        valid_cmp_l4    [1:0]                                                          ; // ���ļ���Ч��־�ȽϽ��

generate
    for (gj = 0; gj < 2; gj = gj + 1) begin: g_pri_cmp_l4
        assign valid_cmp_l4[gj] = valid_cmp_l3[gj*2] | valid_cmp_l3[gj*2+1];
        assign pri_cmp_l4[gj]   = (!valid_cmp_l3[gj*2] && valid_cmp_l3[gj*2+1]) ? pri_cmp_l3[gj*2+1] :
                                  (valid_cmp_l3[gj*2] && !valid_cmp_l3[gj*2+1]) ? pri_cmp_l3[gj*2] :
                                  (valid_cmp_l3[gj*2] && valid_cmp_l3[gj*2+1]) ? 
                                  ((pri_cmp_l3[gj*2] > pri_cmp_l3[gj*2+1]) ? pri_cmp_l3[gj*2] : pri_cmp_l3[gj*2+1]) :
                                  3'b000;
        assign addr_cmp_l4[gj]  = (!valid_cmp_l3[gj*2] && valid_cmp_l3[gj*2+1]) ? addr_cmp_l3[gj*2+1] :
                                  (valid_cmp_l3[gj*2] && !valid_cmp_l3[gj*2+1]) ? addr_cmp_l3[gj*2] :
                                  (valid_cmp_l3[gj*2] && valid_cmp_l3[gj*2+1]) ? 
                                  ((pri_cmp_l3[gj*2] > pri_cmp_l3[gj*2+1]) ? addr_cmp_l3[gj*2] : 
                                   (pri_cmp_l3[gj*2] < pri_cmp_l3[gj*2+1]) ? addr_cmp_l3[gj*2+1] : addr_cmp_l3[gj*2]) :
                                  {QUEUE_ADDR_WIDTH{1'b0}};
    end
endgenerate

// ���弶�Ƚϣ����ձȽ�����
assign r_max_pri   = (!valid_cmp_l4[0] && valid_cmp_l4[1]) ? pri_cmp_l4[1] :
                   (valid_cmp_l4[0] && !valid_cmp_l4[1]) ? pri_cmp_l4[0] :
                   (valid_cmp_l4[0] && valid_cmp_l4[1]) ? 
                   ((pri_cmp_l4[0] > pri_cmp_l4[1]) ? pri_cmp_l4[0] : pri_cmp_l4[1]) :
                   3'b000;

assign r_next_addr = (!valid_cmp_l4[0] && valid_cmp_l4[1]) ? addr_cmp_l4[1] :
                   (valid_cmp_l4[0] && !valid_cmp_l4[1]) ? addr_cmp_l4[0] :
                   (valid_cmp_l4[0] && valid_cmp_l4[1]) ? 
                   ((pri_cmp_l4[0] > pri_cmp_l4[1]) ? addr_cmp_l4[0] : 
                    (pri_cmp_l4[0] < pri_cmp_l4[1]) ? addr_cmp_l4[1] : addr_cmp_l4[0]) :
                   {QUEUE_ADDR_WIDTH{1'b0}};

// ��ǰ�����ַѡ��(�ϸ�������ȼ�)
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_current_process_addr <= {QUEUE_ADDR_WIDTH{1'b0}};
    end else begin
        r_current_process_addr <= ri_cross_metadata_valid_1d == 1'b1 ? r_next_addr : r_current_process_addr;
    end
end

always @(posedge i_clk) begin
    r_process_complete_d1 <= r_process_complete;
end

// ������ɱ�־
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_process_complete <= 1'b0;
    end else begin
        r_process_complete <=   w_is_critical_frame == 1'b1 && o_emac_axi_data_last == 1'd1 ||
                                (w_is_critical_frame == 1'b0) && (((r_timeout_flag == 1'b1) ||
                                ((r_rtag_flag == 1'b1) && (ri_judge_finish == 1'b1) && (ri_discard_en == 1'b1)) ||
                                (w_frame_read_end == 1'd1  && ((r_ack_received & r_ack_expected) == r_ack_expected) && (r_ack_expected != {PORT_NUM{1'b0}}))))
                               ? 1'b1 : 1'b0;
    end
end

/*---------------------------------------- ACK�����߼� -------------------------------------------*/
// ACK���ձ�־����
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_ack_received <= {PORT_NUM{1'b0}};
    end else begin
        r_ack_received <= (ro_mac_cross_axi_data_last == 1'b1) ? {PORT_NUM{1'b0}} :
                          (r_ack_received | ({i_mac_tx7_ack, i_mac_tx6_ack, i_mac_tx5_ack, i_mac_tx4_ack,
                                           i_mac_tx3_ack, i_mac_tx2_ack, i_mac_tx1_ack, i_mac_tx0_ack} & r_ack_expected));
    end
end

// ����ACKͨ��������metadata[59:52]��
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_ack_expected <= {PORT_NUM{1'b0}};
    end else if (ro_tx_req == 1'b1) begin
        r_ack_expected <= w_current_metadata[59:52];
    end
end

/*---------------------------------------- ����������� -------------------------------------------*/
// ����RAM��ָ��
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_data_ram_rd_ptr <= {RAM_ADDR_WIDTH{1'b0}};
    end else begin
        r_data_ram_rd_ptr <=  (w_is_critical_frame == 1'b1 && ri_pass_en == 1'b0 && i_pass_en == 1'b1) || (ro_tx_req == 1'b1) ? r_frame_start_addrs[r_current_process_addr] : 
                              (((r_frame_reading == 1'b1) && (i_mac_cross_axi_data_ready == 1'b1) && 
                               r_frame_end_addr_valid[r_current_process_addr] == 1'b1 && (r_data_ram_rd_ptr == r_frame_end_addrs[r_current_process_addr])) ? r_data_ram_rd_ptr :
                              ((r_frame_reading == 1'b1) && ((i_mac_cross_axi_data_ready == 1'b1) || w_is_critical_frame == 1'b1)) ? (r_data_ram_rd_ptr + {{(RAM_ADDR_WIDTH-1){1'b0}}, 1'b1}) :
                              r_data_ram_rd_ptr);
    end
end

// ֡��ȡ��־
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_frame_reading <= 1'b0;
    end else begin
        r_frame_reading <= (r_current_is_critical == 1'b0 && ro_mac_cross_axi_data_valid == 1'b1 && (r_data_out_cnt >= r_data_out_len - 16'd2) && (i_mac_cross_axi_data_ready == 1'b1)) ? 1'b0 :
                           (r_current_is_critical == 1'b1 && o_emac_axi_data_valid == 1'b1 && (r_data_out_cnt >= r_data_out_len - 16'd1) && (i_emac_axi_data_ready == 1'b1)) ? 1'b0 :
                           (r_current_is_critical == 1'b0 && (r_req_sent == 1'b1) && ((r_ack_received & r_ack_expected) == r_ack_expected) && (r_ack_expected != {PORT_NUM{1'b0}})) ? 1'b1 :
                           (r_current_is_critical == 1'b1 && i_judge_finish == 1'b1 && i_pass_en == 1'd1) ? 1'b1 :
                           r_frame_reading  ;
    end
end

/*---------------------------------------- ��������� -------------------------------------------*/
// �����������ж�last�ź�
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_data_out_cnt <= 16'd0;
    end else begin
        r_data_out_cnt <= (r_current_is_critical == 1'b0 && ro_tx_req == 1'b1) ? 16'd0 :
                          (r_current_is_critical == 1'b1 && r_info_ram_re_d2 == 1'b1) ? 16'd0 :
                          ((ro_mac_cross_axi_data_valid == 1'b1) && (i_mac_cross_axi_data_ready == 1'b1) && r_data_out_cnt <= r_data_out_len) ? (r_data_out_cnt + 16'd1) :
                          ((o_emac_axi_data_valid == 1'b1) && (i_emac_axi_data_ready == 1'b1) && r_data_out_cnt <= r_data_out_len) ? (r_data_out_cnt + 16'd1) :
                          r_data_out_cnt;
    end
end

always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_data_out_len <= 16'd0;
    end else begin
        r_data_out_len <= (r_current_is_critical == 1'b0 && ro_tx_req == 1'b1) ? w_info_ram_rd_data[14:0] : 
                          (r_current_is_critical == 1'b1 && r_info_ram_re_d2 == 1'b1) ? w_info_ram_rd_data[14:0] :
                          r_data_out_len;
    end
end

always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        ro_mac_cross_axi_data_valid <= 1'b0;
    end else begin
        ro_mac_cross_axi_data_valid <= (r_current_is_critical == 1'b0) && (ro_mac_cross_axi_data_valid == 1'd1 && r_data_out_cnt >= r_data_out_len - 1'd1)  ? 1'd0 :
                                     (r_current_is_critical == 1'b0) && ((r_frame_reading == 1'b1) && (r_ack_received != {PORT_NUM{1'b0}})) ? 1'b1 : 1'b0;
    end
end

always @(posedge i_clk) begin
    // ro_mac_cross_axi_data_valid_d1 <= ro_mac_cross_axi_data_valid == 1'd1 && r_data_out_len == r_data_out_cnt ? 1'd0 : ro_mac_cross_axi_data_valid == 1'd1 && r_frame_reading == 1'd1  ? 1'd1 :  1'd0;  
     ro_mac_cross_axi_data_valid_d1 <= ro_mac_cross_axi_data_valid;
end

always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        ro_mac_cross_port_axi_data <= {CROSS_DATA_WIDTH{1'b0}};
    end else begin
        ro_mac_cross_port_axi_data <= (ro_mac_cross_axi_data_valid == 1'b1) ? 
                                      w_data_ram_rd_data[PORT_MNG_DATA_WIDTH + (PORT_MNG_DATA_WIDTH/8)-1:(PORT_MNG_DATA_WIDTH/8)] : 
                                      {CROSS_DATA_WIDTH{1'b0}};
    end
end

always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        ro_mac_cross_axi_data_keep <= {(CROSS_DATA_WIDTH/8){1'b0}};
    end else begin
        ro_mac_cross_axi_data_keep <= (ro_mac_cross_axi_data_valid == 1'b1) ? 
                                      w_data_ram_rd_data[(PORT_MNG_DATA_WIDTH/8)-1:0] : 
                                      {(CROSS_DATA_WIDTH/8){1'b0}};
    end
end

always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        ro_mac_cross_axi_data_last <= 1'b0;
    end else begin
        ro_mac_cross_axi_data_last <= (ro_mac_cross_axi_data_valid == 1'b1 && (r_data_out_cnt == r_data_out_len - 16'd1)) ? 1'b1 : 1'b0;
    end
end

always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        ro_mac_cross_port_axi_user <= 16'b0;
    end else begin
        ro_mac_cross_port_axi_user <= (ro_mac_cross_axi_data_valid == 1'b1) ? w_info_ram_rd_data[15:0] : 16'b0;
    end
end

/*---------------------------------------- ���metadata�� -------------------------------------------*/
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        ro_cross_metadata_valid <= 1'b0;
    end else begin
        ro_cross_metadata_valid <= (r_current_is_critical == 1'b0) && ((ro_tx_req == 1'b1) || (ro_mac_cross_axi_data_valid == 1'd1 && ro_mac_cross_axi_data_valid_d1 == 1'd0))  ? 1'b1 : 1'b0;
    end
end

always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        ro_cross_metadata <= {METADATA_WIDTH{1'b0}};
    end else begin
        ro_cross_metadata <= (r_current_is_critical == 1'b0) && (ro_tx_req == 1'b1) ? w_info_ram_rd_data[FRAME_INFO_WIDTH-1:16] : ro_cross_metadata;
    end
end

always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        ro_cross_metadata_last <= 1'b0;
    end else begin
        ro_cross_metadata_last <= (r_current_is_critical == 1'b0) && ((ro_tx_req == 1'b1) || (ro_mac_cross_axi_data_valid == 1'd1 && ro_mac_cross_axi_data_valid_d1 == 1'd0)) ? 1'b1 : 1'b0;
    end
end

/*---------------------------------------- req����ź� -------------------------------------------*/
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        ro_tx_req <= 1'b0;
    end else begin
        ro_tx_req <= (r_current_is_critical == 1'b0) && (((r_info_ram_re_d2 == 1'd1) && (r_rtag_flag == 1'b0) && (r_queue_empty == 1'b0) && (r_req_sent == 1'b0)) ||
                      ((r_rtag_flag == 1'b1) && (r_cb_result_rcvd == 1'b1) && (r_pass_result == 1'b1) && (r_req_sent == 1'b0))) ? 1'b1 : 1'b0;
    end
end
 

always @(posedge i_clk) begin
    ro_tx_req_d1 <= ro_tx_req;
end 
 
assign w_tx_req = (r_current_is_critical == 1'b0) && ((((r_info_ram_re_d2 == 1'd1) && (r_rtag_flag == 1'b0) && (r_queue_empty == 1'b0) && (r_req_sent == 1'b0)) ||
                  ((r_rtag_flag == 1'b1) && (r_cb_result_rcvd == 1'b1) && (r_pass_result == 1'b1) && (r_req_sent == 1'b0)))) ? 1'b1 : 1'b0;
/*---------------------------------------- �����ֵ -------------------------------------------*/
assign o_mac_axi_data_ready             = ro_mac_axi_data_ready                                            ;
assign o_cross_metadata_ready           = ro_cross_metadata_ready                                          ;
assign o_mac_cross_port_axi_user        = ro_mac_cross_port_axi_user                                       ;
assign o_mac_cross_port_axi_data        = ro_mac_cross_port_axi_data                                       ;
assign o_mac_cross_axi_data_keep        = ro_mac_cross_axi_data_keep                                       ;
// �ؼ�֡��·ʱ������ͨ�������������Ч
assign o_mac_cross_axi_data_valid       = (r_current_is_critical == 1'b1) ? 1'b0 : ro_mac_cross_axi_data_valid_d1 ;
assign o_mac_cross_axi_data_last        = ro_mac_cross_axi_data_last                                       ;
assign o_cross_metadata                 = ro_cross_metadata                                                ;
assign o_cross_metadata_valid           = (r_current_is_critical == 1'b1) ? 1'b0 : ro_cross_metadata_valid      ;
assign o_cross_metadata_last            = ro_cross_metadata_last                                           ;
assign o_rtag_flag                      = ro_rtag_flag                                                     ;
assign o_rtag_squence                   = ro_rtag_squence                                                  ;
assign o_stream_handle                  = ro_stream_handle                                                 ;
assign o_tx_req                         = (r_current_is_critical == 1'b1) ? 1'b0 : ro_tx_req_d1             ;

/*---------------------------------------- �� PORT �ؼ�֡��·��� -------------------------------------------*/   
assign o_emac_port_axi_data    = (r_current_is_critical == 1'b1 && r_frame_reading == 1'b1 && ((r_rtag_flag == 1'b0) || (r_rtag_flag == 1'b1 && r_pass_result == 1'b1))) ? w_data_ram_rd_data[PORT_MNG_DATA_WIDTH + (PORT_MNG_DATA_WIDTH/8)-1:(PORT_MNG_DATA_WIDTH/8)] : {CROSS_DATA_WIDTH{1'b0}};
assign o_emac_port_axi_user    = (r_current_is_critical == 1'b1 && r_frame_reading == 1'b1 && ((r_rtag_flag == 1'b0) || (r_rtag_flag == 1'b1 && r_pass_result == 1'b1))) ? w_info_ram_rd_data[15:0] : 16'b0;
assign o_emac_axi_data_keep    = (r_current_is_critical == 1'b1 && r_frame_reading == 1'b1 && ((r_rtag_flag == 1'b0) || (r_rtag_flag == 1'b1 && r_pass_result == 1'b1))) ? w_data_ram_rd_data[(PORT_MNG_DATA_WIDTH/8)-1:0] : {(CROSS_DATA_WIDTH/8){1'b0}};
assign o_emac_axi_data_valid   = (r_current_is_critical == 1'b1 && r_frame_reading == 1'b1 && ((r_rtag_flag == 1'b0) || (r_rtag_flag == 1'b1 && r_pass_result == 1'b1))) ? 1'b1 : 1'b0;
assign o_emac_axi_data_last    = (r_current_is_critical == 1'b1 && r_frame_reading == 1'b1 && ((r_rtag_flag == 1'b0) || (r_rtag_flag == 1'b1 && r_pass_result == 1'b1)) && (r_data_out_cnt == r_data_out_len - 16'd1)) ? 1'b1 : 1'b0;

assign o_emac_metadata         = (r_current_is_critical == 1'b1 && ((r_rtag_flag == 1'b0) || (r_rtag_flag == 1'b1 && ri_pass_en == 1'b1 && r_pass_result == 1'b1))) ? w_info_ram_rd_data[FRAME_INFO_WIDTH-1:16] : {METADATA_WIDTH{1'b0}};
assign o_emac_metadata_valid   = (r_current_is_critical == 1'b1 && ((r_rtag_flag == 1'b0) || (r_rtag_flag == 1'b1 && ri_pass_en == 1'b1 && r_pass_result == 1'b1))) ? 1'b1 : 1'b0;
assign o_emac_metadata_last    = (r_current_is_critical == 1'b1 && ((r_rtag_flag == 1'b0) || (r_rtag_flag == 1'b1 && ri_pass_en == 1'b1 && r_pass_result == 1'b1))) ? 1'b1 : 1'b0;

/*---------------------------------------- RAM���� -------------------------------------------*/
// ����RAM - �洢֡����
assign w_data_ram_wr_addr = r_data_wr_ptr;
assign w_data_ram_rd_addr = r_data_ram_rd_ptr;
assign w_data_ram_wr_data = {ri_mac_axi_data, ri_mac_axi_data_keep};
assign w_data_ram_we      = (ri_mac_axi_data_valid == 1'b1) && (ro_mac_axi_data_ready == 1'b1);
assign w_data_ram_re      = (r_frame_reading == 1'b1);

ram_simple2port #(
    .RAM_WIDTH               (PORT_MNG_DATA_WIDTH + (PORT_MNG_DATA_WIDTH/8)),
    .RAM_DEPTH               (RAM_DEPTH),
    .RAM_PERFORMANCE         ("LOW_LATENCY"),
    .INIT_FILE               ()
) u_data_ram (
    .addra                   (w_data_ram_wr_addr),
    .addrb                   (w_data_ram_rd_addr),
    .dina                    (w_data_ram_wr_data),
    .clka                    (i_clk),
    .clkb                    (i_clk),
    .wea                     (w_data_ram_we),
    .enb                     (w_data_ram_re),
    .rstb                    (i_rst),
    .regceb                  (1'b1),
    .doutb                   (w_data_ram_rd_data)
);

// ��ϢRAM - �洢֡��Ϣ
assign w_info_ram_wr_addr = r_wr_addr                                                                     ;
assign w_info_ram_rd_addr = r_rd_addr                                                                     ;
assign w_info_ram_wr_data = {ri_cross_metadata, ri_mac_axi_data_user}                                     ;
assign w_info_ram_we      = (ri_cross_metadata_valid == 1'b1) && (ri_cross_metadata_last == 1'b1) && (r_queue_full == 1'b0);

// ��ϢRAM��ʹ�ܣ�ÿ�ν�����һ��ʱ������
// ����������
// 1) r_rd_addr�����仯���л����µĶ����
// 2) �����ɿձ�ǿգ��״���Ч�����ʱ��
reg [QUEUE_ADDR_WIDTH-1:0] r_rd_addr_d1;
reg                        r_queue_empty_d1;
// ���ĵ�ַ�л��ź�
always @(posedge i_clk) begin  
    r_info_ram_we <= w_info_ram_we;
    r_rd_addr_d1 <= r_rd_addr; 
end

// ���Ķ��п��ź�
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_queue_empty_d1 <= 1'b1;
    end else begin
        r_queue_empty_d1 <= r_queue_empty;
    end
end

// ������ϢRAM��ʹ���ź�
always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_info_ram_re <= 1'b0;
    end else begin
        r_info_ram_re <= ((r_rd_addr != r_rd_addr_d1) && r_queue_empty == 1'd0) ? 1'b1 :
                         ((r_queue_empty_d1 == 1'b1) && (r_queue_empty == 1'b0)) ? 1'b1 : 1'b0;
    end
end


always @(posedge i_clk) begin
    if (i_rst == 1'b1) begin
        r_info_ram_re_d1 <= 1'b0;
        r_info_ram_re_d2 <= 1'b0;
    end else begin
        r_info_ram_re_d1 <= r_info_ram_re;
        r_info_ram_re_d2 <= r_info_ram_re_d1;
    end
end


ram_simple2port #(
    .RAM_WIDTH               (FRAME_INFO_WIDTH      ),
    .RAM_DEPTH               (QUEUE_SIZE            ),
    .RAM_PERFORMANCE         ("LOW_LATENCY"         ),
    .INIT_FILE               (                      )
) u_info_ram (
    .addra                   (w_info_ram_wr_addr    ),
    .addrb                   (w_info_ram_rd_addr    ),
    .dina                    (w_info_ram_wr_data    ),
    .clka                    (i_clk                 ),
    .clkb                    (i_clk                 ),
    .wea                     (w_info_ram_we         ),
    .enb                     (r_info_ram_re         ),
    .rstb                    (i_rst                 ),
    .regceb                  (1'b1                  ),
    .doutb                   (w_info_ram_rd_data    )
);

// ��ʱ��״̬�Ĵ��������ֵΪ0
assign o_port_diag_state                = 32'b0;
assign o_port_rx_ultrashort_frm         = 32'b0;
assign o_port_rx_overlength_frm         = 32'b0;
assign o_port_rx_crcerr_frm             = 32'b0;
assign o_port_rx_loopback_frm_cnt       = 32'b0;
assign o_port_broadflow_drop_cnt        = 32'b0;
assign o_port_multiflow_drop_cnt        = 32'b0;
assign o_port_rx_byte_cnt               = 64'b0;
assign o_port_rx_frame_cnt              = 32'b0;
assign o_acl_list_rdy_regs              = 1'b1;

endmodule