/*---------------------------------------- ����ƽ̨�ļܹ� -------------------------------------------*/
`define END_POINTER_SWITCH_CORE
//`define END_POINTER
//`define SWITCH_CORE
/*---------------------------------------- ����CPU��FPGA�����Ľӿ� -----------------------------------*/
`ifdef END_POINTER_SWITCH_CORE
    `define CPU_MAC
    `define MAC1
    `define MAC2
    `define MAC3
    `define MAC4
    `define MAC5
    `define MAC6
    `define MAC7
    `define LLDP
    `define TSN_AS
`elsif END_POINTER
    `define CPU_MAC
    `define MAC1
    `define MAC2
    `define LLDP
    `define TSN_AS
`endif
/*---------------------------------------- ����ƽ̨�ж��ٸ� Mac_port_mng ----------------------------*/

