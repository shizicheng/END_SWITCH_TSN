`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/06/16 09:40:20
// Design Name: 
// Module Name: top_rec
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module qbu_send#(
    parameter                                           AXIS_DATA_WIDTH         =   'd8        ,
    parameter                                           QUEUE_NUM               =   'd8        ,                                                       
    parameter                                           REG_ADDR_BUS_WIDTH      =     8        ,  // ���� MAC ������üĴ�����ַλ��
    parameter                                           REG_DATA_BUS_WIDTH      =     16          // ���� MAC ������üĴ�������λ��
)(
    input           wire                                i_clk                       ,
    input           wire                                i_rst                       ,
    // �Ĵ���д���ƽӿ�     
    //input           wire                                i_switch_reg_bus_we         , // �Ĵ���дʹ��
    //input           wire   [REG_ADDR_BUS_WIDTH-1:0]     i_switch_reg_bus_we_addr    , // �Ĵ���д��ַ
    //input           wire   [REG_DATA_BUS_WIDTH-1:0]     i_switch_reg_bus_we_din     , // �Ĵ���д����
    //input           wire                                i_switch_reg_bus_we_din_v   , // �Ĵ���д����ʹ��
    // �Ĵ��������ƽӿ�     
    //input           wire                                i_switch_reg_bus_rd         , // �Ĵ�����ʹ��
    //input           wire   [REG_ADDR_BUS_WIDTH-1:0]     i_switch_reg_bus_rd_addr    , // �Ĵ�������ַ
    //output          wire   [REG_DATA_BUS_WIDTH-1:0]     o_switch_reg_bus_we_dout    , // �����Ĵ�������
    //output          wire                                o_switch_reg_bus_we_dout_v  , // ��������Чʹ��

    //pmacͨ������
    input           wire    [AXIS_DATA_WIDTH - 1:0]     i_pmac_tx_axis_data         , 
    input           wire    [15:0]                      i_pmac_tx_axis_user         , 
    input           wire    [(AXIS_DATA_WIDTH/8)-1:0]   i_pmac_tx_axis_keep         , 
    input           wire                                i_pmac_tx_axis_last         , 
    input           wire                                i_pmac_tx_axis_valid        , 
    input           wire    [15:0]                      i_pmac_ethertype            , 
    output          wire                                o_pmac_tx_axis_ready        ,
    //emacͨ������
    input           wire    [AXIS_DATA_WIDTH - 1:0]     i_emac_tx_axis_data         , 
    input           wire    [15:0]                      i_emac_tx_axis_user         , 
    input           wire    [(AXIS_DATA_WIDTH/8)-1:0]   i_emac_tx_axis_keep         , 
    input           wire                                i_emac_tx_axis_last         , 
    input           wire                                i_emac_tx_axis_valid        , 
    input           wire    [15:0]                      i_emac_ethertype            ,
    output          wire                                o_emac_tx_axis_ready        ,

    input           wire                                i_qbu_verify_valid          ,
    input           wire                                i_qbu_response_valid        ,

	//
	output			wire								o_send_flag					,
    //������ӿڲ�axi������
    output          wire    [AXIS_DATA_WIDTH - 1:0]     o_mac_axi_data              ,
    output          wire    [(AXIS_DATA_WIDTH/8)-1:0]   o_mac_axi_data_keep         ,
    output          wire                                o_mac_axi_data_valid        ,
    output          wire    [15:0]                      o_mac_axi_data_user         ,
    input           wire                                i_mac_axi_data_ready        ,
    output          wire                                o_mac_axi_data_last         ,
    //ʱ����ź�
    output          wire                                o_mac_time_irq              , // ��ʱ����ж��ź�
    output          wire    [7:0]                       o_mac_frame_seq             , // ֡���к�
    output          wire    [7:0]                       o_timestamp_addr            ,  // ��ʱ����洢�� RAM ��ַ
    //�Ĵ����ӿ�
    output          wire    [7:0]                       o_frag_next_tx              ,
    output          wire                                o_tx_timeout                ,
    output          wire    [15:0]                      o_preempt_success_cnt       ,
    output          wire                                o_preempt_active            ,
    output          wire                                o_preemptable_frame         ,
    output          wire    [15:0]                      o_tx_frames_cnt             ,
    output          wire    [15:0]                      o_tx_fragment_cnt           ,
    output          wire                                o_tx_busy                   ,

    input           wire    [19:0]                      i_watchdog_timer            ,
    input           wire                                i_watchdog_timer_vld        ,
    input           wire    [ 7:0]                      i_min_frag_size             ,
    input           wire                                i_min_frag_size_vld         ,
    input           wire    [ 7:0]                      i_ipg_timer                 ,
    input           wire                                i_ipg_timer_vld             ,

    input           wire                                i_verify_enabled            ,
    input           wire                                i_start_verify              ,
    input           wire                                i_clear_verify              ,
    output 			wire 							    o_verify_succ 		        ,//��֤�ɹ��ź�-
    output 			wire 							    o_verify_succ_val 	        ,//��֤�ɹ���Ч�ź�-
    input           wire    [15:0]                      i_verify_timer		        ,//������֤����֮��ĵȴ�ʱ��
    input  			wire                                i_verify_timer_vld          ,
    output          wire    [15:0]                      o_err_verify_cnt            ,
    output          wire                                o_preempt_enable             //qbu���ܼ���ɹ�
   

    //���������Ҫ���͵�����
    // input           wire    [AXIS_DATA_WIDTH - 1:0]     i_mac_tx_axis_data          ,
    // input           wire    [15:0]                      i_mac_tx_axis_user          , //user�����ݳ�����Ϣ
    // input           wire    [(AXIS_DATA_WIDTH/8)-1:0]   i_mac_tx_axis_keep          , //keep��������
    // input           wire                                i_mac_tx_axis_last          ,
    // input           wire                                i_mac_tx_axis_valid         ,
    // output          wire                                o_mac_tx_axis_ready         ,
    
    // input           wire    [QUEUE_NUM - 1:0]           i_emac_channel_cfg          ,
    // input           wire    [QUEUE_NUM - 1:0]           i_tx_mac_forward_info       , //�ĸ�ͨ���������ݣ��ڲ��趨��Щ���ȼ���eMAC����Щ��pMAC
    // input           wire                                i_tx_mac_forward_info_vld   ,
);            


wire                [AXIS_DATA_WIDTH - 1:0]             o_top_Emac_tx_axis_data  ;  
wire                [15:0]                              o_top_Emac_tx_axis_user  ;  
wire                [(AXIS_DATA_WIDTH/8)-1:0]           o_top_Emac_tx_axis_keep  ;  
wire                                                    o_top_Emac_tx_axis_last  ;  
wire                                                    o_top_Emac_tx_axis_valid ;  
wire                [15:0]                              o_top_Emac_tx_axis_type  ;  

wire                [AXIS_DATA_WIDTH - 1:0]             o_top_Pmac_tx_axis_data  ;
wire                [15:0]                              o_top_Pmac_tx_axis_user  ;
wire                [(AXIS_DATA_WIDTH/8)-1:0]           o_top_Pmac_tx_axis_keep  ;
wire                                                    o_top_Pmac_tx_axis_last  ;
wire                                                    o_top_Pmac_tx_axis_valid ;
wire                [15:0]                              o_top_Pmac_tx_axis_type  ;      

wire                [AXIS_DATA_WIDTH - 1:0]             i_top_Emac_tx_axis_data  ;  
wire                [15:0]                              i_top_Emac_tx_axis_user  ;  
wire                [(AXIS_DATA_WIDTH/8)-1:0]           i_top_Emac_tx_axis_keep  ;  
wire                                                    i_top_Emac_tx_axis_last  ;  
wire                                                    i_top_Emac_tx_axis_valid ;  
wire                [15:0]                              i_top_Emac_tx_axis_type  ;  

wire                [AXIS_DATA_WIDTH - 1:0]             i_top_Pmac_tx_axis_data  ;
wire                [15:0]                              i_top_Pmac_tx_axis_user  ;
wire                [(AXIS_DATA_WIDTH/8)-1:0]           i_top_Pmac_tx_axis_keep  ;
wire                                                    i_top_Pmac_tx_axis_last  ;
wire                                                    i_top_Pmac_tx_axis_valid ;
wire                [15:0]                              i_top_Pmac_tx_axis_type  ;  

//                  FAST_qbu_Emac_tx ��������        
wire                                                    o_emac_send_busy         ;//eamcæ�źţ���ʾemac���ڷ�����
wire                                                    o_emac_send_apply        ;//emac���ݷ�������
wire                                                    i_rx_ready               ;//��֡ģ��׼�������ź�
wire                [15:0]                              o_emac_send_type         ;//Э�����ͣ�����mac֡��ʽ��
wire                [AXIS_DATA_WIDTH-1 :0]              o_emac_send_data         ;//�����ź�
wire                                                    o_emac_send_last         ;//���һ�������ź�
wire                [15:0]                              o_emac_send_len          ;//���ݳ���
wire                                                    o_emac_send_valid        ;//������Ч�ź�
wire                                                    o_emac_smd_val           ;//SMD������Ч�ź�
wire                [15:0]                              o_emac_smd               ;//SMD���� 

//                  mux ��������   
wire    [AXIS_DATA_WIDTH - 1:0]                         i_eth_send_data          ;//�����ź�  
wire    [15:0]                                          i_eth_send_user          ;//������Ϣ  
wire    [(AXIS_DATA_WIDTH/8)-1:0]                       i_eth_send_keep          ;//��������  
wire                                                    i_eth_send_last          ;//���ݽ����ź�
wire                                                    i_eth_send_valid         ;//������Ч�ź� 
wire                                                    o_eth_send_ready         ;//׼���ź�
wire    [15:0]                                          i_eth_send_type          ;//��������
wire                                                    i_eth_smd                ;//SMD����
wire                                                    i_eth_smd_val            ;//SMD������Ч�ź�

wire    [AXIS_DATA_WIDTH - 1:0]                         i_R_rx_axis_data         ;//�����ź�  
wire    [15:0]                                          i_R_rx_axis_user         ;//������Ϣ  
wire    [(AXIS_DATA_WIDTH/8)-1:0]                       i_R_rx_axis_keep         ;//��������  
wire                                                    i_R_rx_axis_last         ;//���ݽ����ź�
//wire                                                  i_R_rx_axis_valid        ;//������Ч�ź�
wire                                                    o_R_rx_axis_ready        ; //׼���ź� 
wire    [AXIS_DATA_WIDTH - 1:0]                         i_V_rx_axis_data         ;//�����ź�  
wire    [15:0]                                          i_V_rx_axis_user         ;//������Ϣ  
wire    [(AXIS_DATA_WIDTH/8)-1:0]                       i_V_rx_axis_keep         ;//��������  
wire                                                    i_V_rx_axis_last         ;//���ݽ����ź�
//wire                                                  i_V_rx_axis_valid        ;//������Ч�ź�
wire                                                    o_V_rx_axis_ready        ; //׼���ź�
                   
wire    [AXIS_DATA_WIDTH - 1:0]                         o_mux_axis_data          ;//�����ź�  
wire    [15:0]                                          o_mux_axis_user          ;//������Ϣ  
wire    [(AXIS_DATA_WIDTH/8)-1:0]                       o_mux_axis_keep          ;//��������  
wire                                                    o_mux_axis_last          ;//���ݽ����ź�
wire                                                    o_mux_axis_valid         ;//������Ч�ź� 
wire                                                    i_mux_axis_ready         ;//׼���ź�
wire    [7:0]                                           o_mux_smd                ;//SMD����
wire                                                    o_mux_smd_val            ;//SMD������Ч�ź�
//wire                                                  o_verify_succ            ;//��֤�ɹ��ź�
//wire                                                  o_verify_succ_val        ;//��֤�ɹ���Ч�ź�
                   
wire                                                    i_pmac_rx_ready          ;//��ģ��׼������
wire    [15:0]                                          o_pmac_send_type         ;//��������
wire    [AXIS_DATA_WIDTH-1 :0]                          o_pmac_send_data         ;//����
wire                                                    o_pmac_send_last         ;//���ݽ����ź�
wire                                                    o_pmac_send_valid        ;//������Ч�ź�
wire    [15:0]                                          o_pmac_send_len          ;//���ݳ���
wire                                                    o_pmac_send_len_val      ;
wire    [15:0]                                          o_pmac_smd               ;//SMD
wire    [15:0]                                          o_pmac_fra               ;//֡������
wire                                                    o_pmac_smd_vld           ;//SMD��Ч�ź�
wire                                                    o_pmac_fra_vld           ;//֡��������Ч�ź�
wire                                                    o_pmac_crc               ;//Ϊ1��Ϊcrc����Ϊmcrc��
                   
wire    [15:0]                                          i_user_set               ;//�û�����(�ݶ����λΪ)
wire                                                    i_user_set_val           ;//�û�������Ч�ź�
wire                                                    i_mac_rx_ready           ;//����֡׼������
wire     [15:0]                                         o_mac_send_type          ;//��������
wire     [AXIS_DATA_WIDTH-1 :0]                         o_mac_send_data          ;//����
wire                                                    o_mac_send_last          ;//���ݽ����ź�
wire    [15:0]                                          o_mac_send_len           ;//���ݳ���
wire                                                    o_mac_send_valid         ;//������Ч�ź�
wire    [15:0]                                          o_mac_smd                ;//SMD
wire    [15:0]                                          o_mac_fra                ;//֡������
wire                                                    o_mac_smd_vld            ;//SMD��Ч�ź�
wire                                                    o_mac_fra_vld            ;//֡��������Ч�ź�
wire                                                    o_mac_crc                ;//Ϊ1��Ϊcrc����Ϊmcrc
wire                                                    o_occupy_succ            ;

wire    [AXIS_DATA_WIDTH - 1:0]     	                o_qbu_verify_data        ;
wire    [15:0]                      	                o_qbu_verify_user        ;
wire    [(AXIS_DATA_WIDTH/8)-1:0]   	                o_qbu_verify_keep        ;
wire                                	                o_qbu_verify_last        ;
wire                                	                o_qbu_verify_valid       ;
wire                                	                i_qbu_verify_ready       ;
wire    [7:0]                       	                o_qbu_verify_smd 	     ;
wire                                                    o_qbu_verify_smd_valid   ;

// wire    [7:0]                                        o_frag_next_tx           ;          
// wire                                                 o_tx_timeout             ;    
// wire    [15:0]                                       o_preempt_success_cnt    ;           
// wire                                                 o_preempt_active         ;    
// wire                                                 o_preemptable_frame      ;
// wire    [15:0]                                       o_tx_frames_cnt          ;
// wire    [15:0]                                       o_tx_fragment_cnt        ; 
// wire                                                 o_tx_busy                ;
                    
// wire    [19:0]                                       i_watchdog_timer         ;    
// wire                                                 i_watchdog_timer_vld     ;
// wire    [ 7:0]                                       i_min_frag_size          ;    
// wire                                                 i_min_frag_size_vld      ;  
// wire    [ 7:0]                                       i_ipg_timer              ;
// wire                                                 i_ipg_timer_vld          ;    

              
// qbu_tx_mac_map #(
//     .AXIS_DATA_WIDTH              (AXIS_DATA_WIDTH),
//     .QUEUE_NUM                    (QUEUE_NUM)
// ) inst_qbu_tx_mac_map (
//     .i_clk                        (i_clk                     ),
//     .i_rst                        (i_rst                     ),
//     .i_mac_tx_axis_data           (i_mac_tx_axis_data        ),
//     .i_mac_tx_axis_keep           (i_mac_tx_axis_keep        ),
//     .i_mac_tx_axis_user           (i_mac_tx_axis_user        ),
//     .i_mac_tx_axis_last           (i_mac_tx_axis_last        ),
//     .i_mac_tx_axis_valid          (i_mac_tx_axis_valid       ),
//     .o_mac_tx_axis_ready          (o_mac_tx_axis_ready       ),

//     .i_emac_channel_cfg           (i_emac_channel_cfg        ),
//     .i_tx_mac_forward_info        (i_tx_mac_forward_info     ),
//     .i_tx_mac_forward_info_vld    (i_tx_mac_forward_info_vld ),
//     .i_verify_succ                (o_verify_succ             ),
//     .i_verify_succ_valid          (o_verify_succ_val         ),

//     .o_emac_tx_axis_data          (i_top_Emac_tx_axis_data   ),
//     .o_emac_tx_axis_user          (i_top_Emac_tx_axis_user   ),
//     .o_emac_tx_axis_keep          (i_top_Emac_tx_axis_keep   ),
//     .o_emac_tx_axis_last          (i_top_Emac_tx_axis_last   ),
//     .o_emac_tx_axis_valid         (i_top_Emac_tx_axis_valid  ),
//     .o_emac_tx_axis_type          (i_top_Emac_tx_axis_type   ),
//     .i_emac_tx_axis_ready         (o_top_Emac_tx_axis_ready  ),

//     .o_pmac_tx_axis_data          (i_top_Pmac_tx_axis_data   ),
//     .o_pmac_tx_axis_user          (i_top_Pmac_tx_axis_user   ),
//     .o_pmac_tx_axis_keep          (i_top_Pmac_tx_axis_keep   ),
//     .o_pmac_tx_axis_last          (i_top_Pmac_tx_axis_last   ),
//     .o_pmac_tx_axis_valid         (i_top_Pmac_tx_axis_valid  ),
//     .o_pmac_tx_axis_type          (i_top_Pmac_tx_axis_type   ),
//     .i_pmac_tx_axis_ready         (o_top_Pmac_tx_axis_ready  )
// );

//��֤��С֡��
    frame_len_detect #(
        .AXIS_DATA_WIDTH                    (AXIS_DATA_WIDTH          )
    ) inst_frame_len_detect (
        .i_clk                              (i_clk                    ),
        .i_rst                              (i_rst                    ),
                    
        .i_top_Emac_tx_axis_data            (i_emac_tx_axis_data      ),
        .i_top_Emac_tx_axis_user            (i_emac_tx_axis_user      ),
        .i_top_Emac_tx_axis_keep            (i_emac_tx_axis_keep      ),
        .i_top_Emac_tx_axis_last            (i_emac_tx_axis_last      ),
        .i_top_Emac_tx_axis_valid           (i_emac_tx_axis_valid     ),
        .i_top_Emac_tx_axis_type            (i_emac_ethertype         ),   
        .o_top_Emac_tx_axis_ready           (o_emac_tx_axis_ready     ),
            
        .i_top_Pmac_tx_axis_data            (i_pmac_tx_axis_data      ),
        .i_top_Pmac_tx_axis_user            (i_pmac_tx_axis_user      ),
        .i_top_Pmac_tx_axis_keep            (i_pmac_tx_axis_keep      ),
        .i_top_Pmac_tx_axis_last            (i_pmac_tx_axis_last      ),
        .i_top_Pmac_tx_axis_valid           (i_pmac_tx_axis_valid     ),
        .i_top_Pmac_tx_axis_type            (i_pmac_ethertype         ),           
        .o_top_Pmac_tx_axis_ready           (o_pmac_tx_axis_ready     ),
            
        .o_top_Emac_tx_axis_data            (o_top_Emac_tx_axis_data  ),
        .o_top_Emac_tx_axis_user            (o_top_Emac_tx_axis_user  ),
        .o_top_Emac_tx_axis_keep            (o_top_Emac_tx_axis_keep  ),
        .o_top_Emac_tx_axis_last            (o_top_Emac_tx_axis_last  ),
        .o_top_Emac_tx_axis_valid           (o_top_Emac_tx_axis_valid ),
        .o_top_Emac_tx_axis_type            (o_top_Emac_tx_axis_type  ),
        .i_top_Emac_tx_axis_ready           (o_top_Emac_tx_axis_ready ),
            
        .o_top_Pmac_tx_axis_data            (o_top_Pmac_tx_axis_data  ),
        .o_top_Pmac_tx_axis_user            (o_top_Pmac_tx_axis_user  ),
        .o_top_Pmac_tx_axis_keep            (o_top_Pmac_tx_axis_keep  ),
        .o_top_Pmac_tx_axis_last            (o_top_Pmac_tx_axis_last  ),
        .o_top_Pmac_tx_axis_valid           (o_top_Pmac_tx_axis_valid ),
        .o_top_Pmac_tx_axis_type            (o_top_Pmac_tx_axis_type  ),
        .i_top_Pmac_tx_axis_ready           (o_top_Pmac_tx_axis_ready )
    );   
    
    qbu_tx_timestamp #(
        .DWIDTH                                 (AXIS_DATA_WIDTH            )
    ) inst_qbu_tx_timestamp(                        
        .i_clk                                  (i_clk                      ),
        .i_rst                                  (i_rst                      ),
        .i_mac_axis_data                        (o_mac_axi_data             ),
        .i_mac_axis_valid                       (o_mac_axi_data_valid       ),
        .o_mac_time_irq                         (o_mac_time_irq             ), // ��Ҫ���ӻ�����
        .o_mac_frame_seq                        (o_mac_frame_seq            ), // ��Ҫ���ӻ�����
        .o_timestamp_addr                       (o_timestamp_addr           )  // ��Ҫ���ӻ�����
    );

    FAST_qbu_Emac_tx    #(
        .AXIS_DATA_WIDTH                        (AXIS_DATA_WIDTH            )
    ) inst_FAST_qbu_Emac_tx    (    
        .i_clk                                  (i_clk                      ),   
        .i_rst                                  (i_rst                      ),
        //����emacͨ������׼������  
        .i_top_Emac_tx_axis_data                (o_top_Emac_tx_axis_data    ),   
        .i_top_Emac_tx_axis_user                (o_top_Emac_tx_axis_user    ),   
        .i_top_Emac_tx_axis_keep                (o_top_Emac_tx_axis_keep    ),   
        .i_top_Emac_tx_axis_last                (o_top_Emac_tx_axis_last    ),   
        .i_top_Emac_tx_axis_valid               (o_top_Emac_tx_axis_valid   ),   
        .i_top_Emac_tx_axis_type                (o_top_Emac_tx_axis_type    ),   
        .o_top_Emac_tx_axis_ready               (o_top_Emac_tx_axis_ready   ),
        //�����Muxģ�� 
        .i_pmac_send_busy                       (o_pamc_send_busy           ),
        .i_pmac_send_apply                      (o_pamc_send_apply          ),
        .o_emac_send_busy                       (o_emac_send_busy           ),
        .o_emac_send_apply                      (o_emac_send_apply          ),
        .i_rx_ready                             (o_emac_rx_ready            ),
        .o_emac_data_noempty                    (o_emac_data_noempty        ),
        .o_send_type                            (o_emac_send_type           ),
        .o_send_data                            (o_emac_send_data           ),
        .o_send_last                            (o_emac_send_last           ),
        .o_send_valid                           (o_emac_send_valid          ),
        .o_smd_val                              (o_emac_smd_val             ),
        .o_send_len                             (o_emac_send_len            ),
        .o_smd                                  (o_emac_smd                 )                  
    );

    Mux #(
      .AXIS_DATA_WIDTH  (AXIS_DATA_WIDTH)
    ) inst_Mux    (
        .i_clk                                  (i_clk                      ),   
        .i_rst                                  (i_rst                      ),

        .i_eth_send_data                        (i_eth_send_data            ),
        .i_eth_send_user                        (i_eth_send_user            ),
        .i_eth_send_keep                        (i_eth_send_keep            ),
        .i_eth_send_last                        (i_eth_send_last            ),
        .i_eth_send_valid                       (i_eth_send_valid           ),
        .o_eth_send_ready                       (o_eth_send_ready           ),
        .i_eth_send_type                        (i_eth_send_type            ),
        .i_eth_smd                              (i_eth_smd                  ),
        .i_eth_smd_val                          (i_eth_smd_val              ),

        .i_verify_send_data                     (o_qbu_verify_data          ),
        .i_verify_send_user                     (o_qbu_verify_user          ),
        .i_verify_send_keep                     (o_qbu_verify_keep          ),
        .i_verify_send_last                     (o_qbu_verify_last          ),
        .i_verify_send_valid                    (o_qbu_verify_valid         ),
        .o_verify_send_ready                    (i_qbu_verify_ready         ),
        .i_verify_smd                           (o_qbu_verify_smd           ),
        .i_verify_smd_val                       (o_qbu_verify_smd_valid     ),

        .i_verify_succ                          (o_verify_succ              ),
        .i_verify_succ_val                      (o_verify_succ_val          ),

        .o_pmac_rx_ready                        (i_pmac_rx_ready            ),
        .i_pmac_send_type                       (o_pmac_send_type           ),
        .i_pmac_send_data                       (o_pmac_send_data           ),
        .i_pmac_send_last                       (o_pmac_send_last           ),
        .i_pmac_send_valid                      (o_pmac_send_valid          ),
        .i_pmac_send_len                        (o_pmac_send_len            ),
        .i_pmac_smd                             (o_pmac_smd                 ),
        .i_pmac_fra                             (o_pmac_fra                 ),
        .i_pmac_smd_vld                         (o_pmac_smd_vld             ),
        .i_pmac_fra_vld                         (o_pmac_fra_vld             ),
        .i_pmac_crc                             (o_pmac_crc                 ),

        .o_emac_rx_ready                        (o_emac_rx_ready            ),
        .i_emac_send_type                       (o_emac_send_type           ),
        .i_emac_send_data                       (o_emac_send_data           ),
        .i_emac_send_len                        (o_emac_send_len            ),
        .i_emac_send_last                       (o_emac_send_last           ),
        .i_emac_send_valid                      (o_emac_send_valid          ),
        .i_emac_smd_val                         (o_emac_smd_val             ),
        .i_emac_smd                             (o_emac_smd                 ),
        // 
        .i_mac_rx_ready                         (o_udp_ready                ),
        .o_mac_send_type                        (o_mac_send_type            ),
        .o_mac_send_data                        (o_mac_send_data            ),
        .o_mac_send_last                        (o_mac_send_last            ),
        .o_mac_send_valid                       (o_mac_send_valid           ),
        .o_mac_send_len                         (o_mac_send_len             ),
        .o_mac_smd                              (o_mac_smd                  ),
        .o_mac_fra                              (o_mac_fra                  ),
        .o_mac_smd_vld                          (o_mac_smd_vld              ),
        .o_mac_fra_vld                          (o_mac_fra_vld              ),
        .o_mac_crc                              (o_mac_crc                  )  
    );

    MAC_tx #(
      .AXIS_DATA_WIDTH  (AXIS_DATA_WIDTH)
    ) inst_MAC_tx    (
        .i_clk                                  (i_clk                      ),   
        .i_rst                                  (i_rst                      ),
        .i_target_mac                           (i_target_mac               ),
        .i_target_mac_valid                     (i_target_mac_valid         ),
        .i_source_mac                           (i_source_mac               ),
        .i_source_mac_valid                     (i_source_mac_valid         ),
        .o_udp_ready                            (o_udp_ready                ),

        .i_send_type                            (o_mac_send_type            ),
        .i_send_len                             (o_mac_send_len             ),
        .i_pmac_send_len_val                    (o_pmac_send_len_val        ),
        .i_pmac_send_len                        (o_pmac_send_len            ),
        .i_send_data                            (o_mac_send_data            ),
        .i_send_last                            (o_mac_send_last            ),
        .i_send_valid                           (o_mac_send_valid           ),
        .i_smd                                  (o_mac_smd                  ),
        .i_fra                                  (o_mac_fra                  ),
        .i_smd_vld                              (o_mac_smd_vld              ),
        .i_fra_vld                              (o_mac_fra_vld              ),
        .i_crc                                  (o_mac_crc                  ),
        .i_eamc_send_busy                       (o_emac_send_busy           ),
        .i_pamc_send_busy                       (o_emac_send_apply          ),
		//
		.o_send_flag							(o_send_flag				),
        //�����phy�ӿڲ�
        .o_mac_axi_data                         (o_mac_axi_data             ),  
        .o_mac_axi_data_keep                    (o_mac_axi_data_keep        ),  
        .o_mac_axi_data_valid                   (o_mac_axi_data_valid       ),  
        .o_mac_axi_data_user                    (o_mac_axi_data_user        ),  
        .i_mac_axi_data_ready                   (i_mac_axi_data_ready       ),  
        .o_mac_axi_data_last                    (o_mac_axi_data_last        ),  
        //�Ĵ����ӿ�    
        .o_tx_frames_cnt                        (o_tx_frames_cnt            ),    
        .o_tx_fragment_cnt                      (o_tx_fragment_cnt          ),    
        .i_ipg_timer                            (i_ipg_timer                ),    
        .i_ipg_timer_vld                        (i_ipg_timer_vld            ),    
        .o_tx_busy                              (o_tx_busy                  )   
    );

    FAST_qbu_Pmac_tx  #(
        .AXIS_DATA_WIDTH  (AXIS_DATA_WIDTH)
    )inst_FAST_qbu_Pmac_tx(
        .i_clk                                  ( i_clk                       ),
        .i_rst                                  ( i_rst                       ),
        .i_top_Pmac_tx_axis_data                (o_top_Pmac_tx_axis_data      ),
        .i_top_Pmac_tx_axis_user                (o_top_Pmac_tx_axis_user      ),
        .i_top_Pmac_tx_axis_keep                (o_top_Pmac_tx_axis_keep      ),
        .i_top_Pmac_tx_axis_last                (o_top_Pmac_tx_axis_last      ),
        .i_top_Pmac_tx_axis_valid               (o_top_Pmac_tx_axis_valid     ),
        .i_top_Pmac_tx_axis_type                (o_top_Pmac_tx_axis_type      ),
        .o_pmac_send_len                        (o_pmac_send_len              ),
        .o_pmac_send_len_val                    (o_pmac_send_len_val          ),
        .i_emac_send_busy                       (o_emac_send_busy             ),
        .i_emac_data_noempty                    (o_emac_data_noempty          ),
        .i_emac_send_apply                      (o_emac_send_apply            ),
        .i_rx_ready                             (i_pmac_rx_ready              ),
        .o_top_Pmac_tx_axis_ready               (o_top_Pmac_tx_axis_ready     ),
        .o_pamc_send_busy                       (o_pamc_send_busy             ),
        .o_pamc_send_apply                      (o_pamc_send_apply            ),
        .o_send_type                            (o_pmac_send_type             ),
        .o_send_data                            (o_pmac_send_data             ),
        .o_send_last                            (o_pmac_send_last             ),
        .o_send_valid                           (o_pmac_send_valid            ),
        .o_smd                                  (o_pmac_smd                   ),
        .o_fra                                  (o_pmac_fra                   ),
        .o_smd_vld                              (o_pmac_smd_vld               ),
        .o_fra_vld                              (o_pmac_fra_vld               ),
        .o_crc                                  (o_pmac_crc                   ),
        //�Ĵ����ӿ�                    
        .o_frag_next_tx                         (o_frag_next_tx               ),     
        .i_watchdog_timer                       (i_watchdog_timer             ),     
        .i_watchdog_timer_vld                   (i_watchdog_timer_vld         ),     
        .o_tx_timeout                           (o_tx_timeout                 ),     
        .o_preempt_success_cnt                  (o_preempt_success_cnt        ),     
        .i_min_frag_size                        (i_min_frag_size              ),     
        .i_min_frag_size_vld                    (i_min_frag_size_vld          ),     
        .o_preempt_active                       (o_preempt_active             ),     
        .o_preemptable_frame                    (o_preemptable_frame          )   
    );

    verified #(
        .AXIS_DATA_WIDTH                        (AXIS_DATA_WIDTH            )
    ) inst_verified (                             
        .i_clk                                  (i_clk                      ),
        .i_rst                                  (i_rst                      ),

        .i_qbu_verify_valid                     (i_qbu_verify_valid         ),
        .i_qbu_response_valid                   (i_qbu_response_valid       ),
        
        .o_verify_succ                          (o_verify_succ              ),
        .o_verify_succ_val                      (o_verify_succ_val          ),
        // verified_to_txmac
        .o_qbu_verify_data                      (o_qbu_verify_data          ), 
        .o_qbu_verify_user                      (o_qbu_verify_user          ), 
        .o_qbu_verify_keep                      (o_qbu_verify_keep          ), 
        .o_qbu_verify_last                      (o_qbu_verify_last          ), 
        .o_qbu_verify_valid                     (o_qbu_verify_valid         ), 
        .i_qbu_verify_ready                     (i_qbu_verify_ready         ), 
        .o_qbu_verify_smd                       (o_qbu_verify_smd           ), 
        .o_qbu_verify_smd_valid                 (o_qbu_verify_smd_valid     ), 
        //�Ĵ����ź�
        .i_verify_enabled                       (i_verify_enabled           ),
        .i_start_verify                         (i_start_verify             ),
        .i_clear_verify                         (i_clear_verify             ),
        .i_verify_timer                         (i_verify_timer             ),
        .i_verify_timer_vld                     (i_verify_timer_vld         ),
        .o_err_verify_cnt                       (o_err_verify_cnt           ),
        .o_preempt_enable                       (o_preempt_enable           )
    );
/*
    qbu_tx_reg inst_qbu_tx_reg (
        .i_clk                      (i_clk                      ),
        .i_rst                      (i_rst                      ),
        // .i_qbu_bus_we           (i_qbu_bus_we               ),
        // .i_qbu_bus_addr         (i_qbu_bus_addr             ),
        // .i_qbu_bus_din          (i_qbu_bus_din              ),
        // .i_qbu_bus_rd           (i_qbu_bus_rd               ),
        .i_switch_reg_bus_we        (i_switch_reg_bus_we       ),
        .i_switch_reg_bus_we_addr   (i_switch_reg_bus_we_addr  ),
        .i_switch_reg_bus_we_din    (i_switch_reg_bus_we_din   ),
        .i_switch_reg_bus_we_din_v  (i_switch_reg_bus_we_din_v ),
        .i_switch_reg_bus_rd        (i_switch_reg_bus_rd       ),
        .i_switch_reg_bus_rd_addr   (i_switch_reg_bus_rd_addr  ),
        .o_switch_reg_bus_we_dout   (o_switch_reg_bus_we_dout  ),
        .o_switch_reg_bus_we_dout_v (o_switch_reg_bus_we_dout_v),

        .i_tx_busy                  (o_tx_busy                  ),
        .i_preemptable_frame        (o_preemptable_frame        ),
        .i_preempt_active           (o_preempt_active           ),
        .i_preempt_enable           (o_preempt_enable           ),
        .i_tx_fragment_cnt          (o_tx_fragment_cnt          ),
        .i_err_verify_cnt           (o_err_verify_cnt           ),
        .i_tx_frames_cnt            (o_tx_frames_cnt            ),
        .i_preempt_success_cnt      (o_preempt_success_cnt      ),
        .i_tx_timeout               (o_tx_timeout               ),
        .i_frag_next_tx             (o_frag_next_tx             ),

        .o_verify_enabled           (i_verify_enabled           ),
        .o_min_frag_size            (i_min_frag_size            ),
        .o_min_frag_size_valid      (i_min_frag_size_vld        ),
        .o_verify_timer             (i_verify_timer             ),
        .o_verify_timer_valid       (i_verify_timer_vld         ),
        .o_ipg_timer                (i_ipg_timer                ),
        .o_ipg_timer_valid          (i_ipg_timer_vld            ),
        .o_reset                    (o_reset                    ),
        .o_start_verify             (i_start_verify             ),
        .o_clear_verify             (i_clear_verify             ),
        .o_watchdog_timer           (i_watchdog_timer           ),
        .o_watchdog_timer_valid     (i_watchdog_timer_vld       ) 

        // .o_qbu_bus_dout             (o_qbu_bus_dout             )
    );
*/
/*
    ila_0 your_inst_ila_0 (
    .i_clk(i_clk), // input wire i_clk


    .probe0(o_pmac_send_data        ), // input wire [7:0]  probe0  
    .probe1(o_pmac_send_valid   ), // input wire [0:0]  probe1 
    .probe2(o_emac_send_data        ), // input wire [7:0]  probe2 
    .probe3(o_emac_send_valid   )
);
*/
endmodule
