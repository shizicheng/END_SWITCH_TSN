`define CPU_MAC
`define MAC1
`define MAC2
`define MAC3
`define MAC4
`define MAC5
`define MAC6
`define MAC7
module rx_mac_reg#(
    parameter                                                   PORT_NUM                =      8        ,  // �������Ķ˿���
    parameter                                                   REG_ADDR_BUS_WIDTH      =      8        ,  // ���� MAC ������üĴ�����ַλ��
    parameter                                                   REG_DATA_BUS_WIDTH      =      32         // ���� MAC ������üĴ�������λ��
)(
    input               wire                                    i_clk                               ,   // 250MHz
    input               wire                                    i_rst                               ,
    /*---------------------------------------- ƽ̨�Ĵ��������� RXMAC ��صļĴ��� -------------------------------------------*/
`ifdef CPU_MAC
    output              wire   [15:0]                           o_hash_ploy_regs_0                  , // ��ϣ����ʽ
    output              wire   [15:0]                           o_hash_init_val_regs_0              , // ��ϣ����ʽ��ʼֵ
    output              wire                                    o_hash_regs_vld_0                   ,
    output              wire                                    o_port_rxmac_down_regs_0            , // �˿ڽ��շ���MAC�ر�ʹ��
    output              wire                                    o_port_broadcast_drop_regs_0        , // �˿ڹ㲥֡����ʹ��
    output              wire                                    o_port_multicast_drop_regs_0        , // �˿��鲥֡����ʹ��
    output              wire                                    o_port_loopback_drop_regs_0         , // �˿ڻ���֡����ʹ��
    output              wire   [47:0]                           o_port_mac_regs_0                   , // �˿ڵ� MAC ��ַ
    output              wire                                    o_port_mac_vld_regs_0               , // ʹ�ܶ˿� MAC ��ַ��Ч
    output              wire   [7:0]                            o_port_mtu_regs_0                   , // MTU����ֵ
    output              wire   [PORT_NUM-1:0]                   o_port_mirror_frwd_regs_0           , // ����ת���Ĵ���������Ӧ�Ķ˿���1���򱾶˿ڽ��յ����κ�ת������֡������ת��ֵ����1�Ķ˿�
    output              wire   [15:0]                           o_port_flowctrl_cfg_regs_0          , // ������������
    output              wire   [4:0]                            o_port_rx_ultrashortinterval_num_0  , // ֡���
    // ACL �Ĵ���
    output              wire   [PORT_NUM-1:0]                   o_acl_port_sel_0                     , // ѡ��Ҫ���õĶ˿�
    output              wire                                    o_acl_clr_list_regs_0                , // ��ռĴ����б�
    input               wire                                    i_acl_list_rdy_regs_0                , // ���üĴ�����������
    output              wire   [4:0]                            o_acl_item_sel_regs_0                , // ������Ŀѡ��
    //output              wire   [5:0]                            o_acl_item_waddr_regs_0              , // ÿ����Ŀ���֧�ֱȶ� 64 �ֽ�
    //output              wire   [7:0]                            o_acl_item_din_regs_0                , // ��Ҫ�Ƚϵ��ֽ�����
    //output              wire                                    o_acl_item_we_regs_0                 , // ����ʹ���ź�
    //output              wire   [15:0]                           o_acl_item_rslt_regs_0               , // ƥ��Ľ��ֵ - [7:0] ���֡����, [15:8] ACLת��ָ���˿�
    //output              wire                                    o_acl_item_complete_regs_0           , // �˿� ACL �����������ʹ���ź�
    output              wire   [95:0]                           o_acl_item_dmac_code_0                ,
    output              wire   [95:0]                           o_acl_item_smac_code_0                ,
    output              wire   [63:0]                           o_acl_item_vlan_code_0                ,
    output              wire   [31:0]                           o_acl_item_ethtype_code_0             ,
    output              wire   [5:0]                            o_acl_item_action_pass_state_0        ,
    output              wire   [15:0]                           o_acl_item_action_cb_streamhandle_0   ,
    output              wire   [5:0]                            o_acl_item_action_flowctrl_0          ,
    output              wire   [15:0]                           o_acl_item_action_txport_0            ,
    // ״̬�Ĵ���
    input              wire   [15:0]                            i_port_diag_state_0                  , // �˿�״̬�Ĵ�����������Ĵ�����˵������ 
    // ��ϼĴ���
    input              wire                                     i_port_rx_ultrashort_frm_0           , // �˿ڽ��ճ���֡(С��64�ֽ�)
    input              wire                                     i_port_rx_overlength_frm_0           , // �˿ڽ��ճ���֡(����MTU�ֽ�)
    input              wire                                     i_port_rx_crcerr_frm_0               , // �˿ڽ���CRC����֡
    input              wire  [15:0]                             i_port_rx_loopback_frm_cnt_0         , // �˿ڽ��ջ���֡������ֵ
    input              wire  [15:0]                             i_port_broadflow_drop_cnt_0          , // �˿ڽ��յ��㲥������������֡������ֵ
    input              wire  [15:0]                             i_port_multiflow_drop_cnt_0          , // �˿ڽ��յ��鲥������������֡������ֵ
    // ����ͳ�ƼĴ���
    input              wire  [15:0]                             i_port_rx_byte_cnt_0                 , // �˿�0�����ֽڸ���������ֵ
    input              wire  [15:0]                             i_port_rx_frame_cnt_0                ,  // �˿�0����֡����������ֵ  

    //qbu_rx�Ĵ���  
    input              wire                                     i_rx_busy_0                          , // ����æ�ź�
    input              wire  [15:0]                             i_rx_fragment_cnt_0                  , // ���շ�Ƭ����
    input              wire                                     i_rx_fragment_mismatch_0             , // ��Ƭ��ƥ��
    input              wire  [15:0]                             i_err_rx_crc_cnt_0                   , // CRC�������
    input              wire  [15:0]                             i_err_rx_frame_cnt_0                 , // ֡�������
    input              wire  [15:0]                             i_err_fragment_cnt_0                 , // ��Ƭ�������
    input              wire  [15:0]                             i_rx_frames_cnt_0                    , // ����֡����
    input              wire  [7:0]                              i_frag_next_rx_0                     , // ��һ����Ƭ��
    input              wire  [7:0]                              i_frame_seq_0                        , // ֡���
    output             wire                                     o_reset_0                            ,
`endif
`ifdef MAC1
    output              wire   [15:0]                           o_hash_ploy_regs_1                  , // ��ϣ����ʽ
    output              wire   [15:0]                           o_hash_init_val_regs_1              , // ��ϣ����ʽ��ʼֵ
    output              wire                                    o_hash_regs_vld_1                   ,
    output              wire                                    o_port_rxmac_down_regs_1            , // �˿ڽ��շ���MAC�ر�ʹ��
    output              wire                                    o_port_broadcast_drop_regs_1        , // �˿ڹ㲥֡����ʹ��
    output              wire                                    o_port_multicast_drop_regs_1        , // �˿��鲥֡����ʹ��
    output              wire                                    o_port_loopback_drop_regs_1         , // �˿ڻ���֡����ʹ��
    output              wire   [47:0]                           o_port_mac_regs_1                   , // �˿ڵ� MAC ��ַ
    output              wire                                    o_port_mac_vld_regs_1               , // ʹ�ܶ˿� MAC ��ַ��Ч
    output              wire   [7:0]                            o_port_mtu_regs_1                   , // MTU����ֵ
    output              wire   [PORT_NUM-1:0]                   o_port_mirror_frwd_regs_1           , // ����ת���Ĵ���������Ӧ�Ķ˿���1���򱾶˿ڽ��յ����κ�ת������֡������ת��ֵ����1�Ķ˿�
    output              wire   [15:0]                           o_port_flowctrl_cfg_regs_1          , // ������������
    output              wire   [4:0]                            o_port_rx_ultrashortinterval_num_1  , // ֡���
    // ACL �Ĵ�
    output              wire   [PORT_NUM-1:0]                   o_acl_port_sel_1                     , // ѡ��Ҫ���õĶ˿�
    output              wire                                    o_acl_clr_list_regs_1                , // ��ռĴ����б�
    input               wire                                    i_acl_list_rdy_regs_1                , // ���üĴ�����������
    output              wire   [4:0]                            o_acl_item_sel_regs_1                , // ������Ŀѡ��
    //output              wire   [5:0]                            o_acl_item_waddr_regs_1              , // ÿ����Ŀ���֧�ֱȶ� 64 �ֽ�
    //output              wire   [7:0]                            o_acl_item_din_regs_1                , // ��Ҫ�Ƚϵ��ֽ�����
    //output              wire                                    o_acl_item_we_regs_1                 , // ����ʹ���ź�
    //output              wire   [15:0]                           o_acl_item_rslt_regs_1               , // ƥ��Ľ��ֵ - [7:0] ���֡����, [15:8] ACLת��ָ���˿�
    //output              wire                                    o_acl_item_complete_regs_1           , // �˿� ACL �����������ʹ���ź�
    output              wire   [95:0]                           o_acl_item_dmac_code_1                ,
    output              wire   [95:0]                           o_acl_item_smac_code_1                ,
    output              wire   [63:0]                           o_acl_item_vlan_code_1                ,
    output              wire   [31:0]                           o_acl_item_ethtype_code_1             ,
    output              wire   [5:0]                            o_acl_item_action_pass_state_1        ,
    output              wire   [15:0]                           o_acl_item_action_cb_streamhandle_1   ,
    output              wire   [5:0]                            o_acl_item_action_flowctrl_1          ,
    output              wire   [15:0]                           o_acl_item_action_txport_1            ,
    // ״̬�Ĵ���
    input              wire   [15:0]                            i_port_diag_state_1                  , // �˿�״̬�Ĵ�����������Ĵ�����˵������ 
    // ��ϼĴ���
    input              wire                                     i_port_rx_ultrashort_frm_1           , // �˿ڽ��ճ���֡(С��64�ֽ�)
    input              wire                                     i_port_rx_overlength_frm_1           , // �˿ڽ��ճ���֡(����MTU�ֽ�)
    input              wire                                     i_port_rx_crcerr_frm_1               , // �˿ڽ���CRC����֡
    input              wire  [15:0]                             i_port_rx_loopback_frm_cnt_1         , // �˿ڽ��ջ���֡������ֵ
    input              wire  [15:0]                             i_port_broadflow_drop_cnt_1          , // �˿ڽ��յ��㲥������������֡������ֵ
    input              wire  [15:0]                             i_port_multiflow_drop_cnt_1          , // �˿ڽ��յ��鲥������������֡������ֵ
    // ����ͳ�ƼĴ���
    input              wire  [15:0]                             i_port_rx_byte_cnt_1                 , // �˿�0�����ֽڸ���������ֵ
    input              wire  [15:0]                             i_port_rx_frame_cnt_1                , // �˿�0����֡����������ֵ  

    //qbu_rx�Ĵ���  
    input              wire                                     i_rx_busy_1                          , // ����æ�ź�
    input              wire  [15:0]                             i_rx_fragment_cnt_1                  , // ���շ�Ƭ����
    input              wire                                     i_rx_fragment_mismatch_1             , // ��Ƭ��ƥ��
    input              wire  [15:0]                             i_err_rx_crc_cnt_1                   , // CRC�������
    input              wire  [15:0]                             i_err_rx_frame_cnt_1                 , // ֡�������
    input              wire  [15:0]                             i_err_fragment_cnt_1                 , // ��Ƭ�������
    input              wire  [15:0]                             i_rx_frames_cnt_1                    , // ����֡����
    input              wire  [7:0]                              i_frag_next_rx_1                     , // ��һ����Ƭ��
    input              wire  [7:0]                              i_frame_seq_1                        , // ֡���
    output             wire                                     o_reset_1                            ,
`endif
`ifdef MAC2
    output              wire   [15:0]                           o_hash_ploy_regs_2                  , // ��ϣ����ʽ
    output              wire   [15:0]                           o_hash_init_val_regs_2              , // ��ϣ����ʽ��ʼֵ
    output              wire                                    o_hash_regs_vld_2                   ,
    output              wire                                    o_port_rxmac_down_regs_2            , // �˿ڽ��շ���MAC�ر�ʹ��
    output              wire                                    o_port_broadcast_drop_regs_2        , // �˿ڹ㲥֡����ʹ��
    output              wire                                    o_port_multicast_drop_regs_2        , // �˿��鲥֡����ʹ��
    output              wire                                    o_port_loopback_drop_regs_2         , // �˿ڻ���֡����ʹ��
    output              wire   [47:0]                           o_port_mac_regs_2                   , // �˿ڵ� MAC ��ַ
    output              wire                                    o_port_mac_vld_regs_2               , // ʹ�ܶ˿� MAC ��ַ��Ч
    output              wire   [7:0]                            o_port_mtu_regs_2                   , // MTU����ֵ
    output              wire   [PORT_NUM-1:0]                   o_port_mirror_frwd_regs_2           , // ����ת���Ĵ���������Ӧ�Ķ˿���1���򱾶˿ڽ��յ����κ�ת������֡������ת��ֵ����1�Ķ˿�
    output              wire   [15:0]                           o_port_flowctrl_cfg_regs_2          , // ������������
    output              wire   [4:0]                            o_port_rx_ultrashortinterval_num_2  , // ֡���
    // ACL �Ĵ�
    output              wire   [PORT_NUM-1:0]                   o_acl_port_sel_2                     , // ѡ��Ҫ���õĶ˿�
    output              wire                                    o_acl_clr_list_regs_2                , // ��ռĴ����б�
    input               wire                                    i_acl_list_rdy_regs_2                , // ���üĴ�����������
    output              wire   [4:0]                            o_acl_item_sel_regs_2                , // ������Ŀѡ��
    //output              wire   [5:0]                            o_acl_item_waddr_regs_2              , // ÿ����Ŀ���֧�ֱȶ� 64 �ֽ�
    //output              wire   [7:0]                            o_acl_item_din_regs_2                , // ��Ҫ�Ƚϵ��ֽ�����
    //output              wire                                    o_acl_item_we_regs_2                 , // ����ʹ���ź�
    //output              wire   [15:0]                           o_acl_item_rslt_regs_2               , // ƥ��Ľ��ֵ - [7:0] ���֡����, [15:8] ACLת��ָ���˿�
    //output              wire                                    o_acl_item_complete_regs_2           , // �˿� ACL �����������ʹ���ź�
    output              wire   [95:0]                           o_acl_item_dmac_code_2                ,
    output              wire   [95:0]                           o_acl_item_smac_code_2                ,
    output              wire   [63:0]                           o_acl_item_vlan_code_2                ,
    output              wire   [31:0]                           o_acl_item_ethtype_code_2             ,
    output              wire   [5:0]                            o_acl_item_action_pass_state_2        ,
    output              wire   [15:0]                           o_acl_item_action_cb_streamhandle_2   ,
    output              wire   [5:0]                            o_acl_item_action_flowctrl_2          ,
    output              wire   [15:0]                           o_acl_item_action_txport_2            ,
    // ״̬�Ĵ���
    input              wire   [15:0]                            i_port_diag_state_2                  , // �˿�״̬�Ĵ�����������Ĵ�����˵������ 
    // ��ϼĴ���
    input              wire                                     i_port_rx_ultrashort_frm_2           , // �˿ڽ��ճ���֡(С��64�ֽ�)
    input              wire                                     i_port_rx_overlength_frm_2           , // �˿ڽ��ճ���֡(����MTU�ֽ�)
    input              wire                                     i_port_rx_crcerr_frm_2               , // �˿ڽ���CRC����֡
    input              wire  [15:0]                             i_port_rx_loopback_frm_cnt_2         , // �˿ڽ��ջ���֡������ֵ
    input              wire  [15:0]                             i_port_broadflow_drop_cnt_2          , // �˿ڽ��յ��㲥������������֡������ֵ
    input              wire  [15:0]                             i_port_multiflow_drop_cnt_2          , // �˿ڽ��յ��鲥������������֡������ֵ
    // ����ͳ�ƼĴ���
    input              wire  [15:0]                             i_port_rx_byte_cnt_2                 , // �˿�0�����ֽڸ���������ֵ
    input              wire  [15:0]                             i_port_rx_frame_cnt_2                ,  // �˿�0����֡����������ֵ 

    //qbu_rx�Ĵ���  
    input              wire                                     i_rx_busy_2                          , // ����æ�ź�
    input              wire  [15:0]                             i_rx_fragment_cnt_2                  , // ���շ�Ƭ����
    input              wire                                     i_rx_fragment_mismatch_2             , // ��Ƭ��ƥ��
    input              wire  [15:0]                             i_err_rx_crc_cnt_2                   , // CRC�������
    input              wire  [15:0]                             i_err_rx_frame_cnt_2                 , // ֡�������
    input              wire  [15:0]                             i_err_fragment_cnt_2                 , // ��Ƭ�������
    input              wire  [15:0]                             i_rx_frames_cnt_2                    , // ����֡����
    input              wire  [7:0]                              i_frag_next_rx_2                     , // ��һ����Ƭ��
    input              wire  [7:0]                              i_frame_seq_2                        , // ֡���
    output             wire                                     o_reset_2                            ,
`endif
`ifdef MAC3
    output              wire   [15:0]                           o_hash_ploy_regs_3                 , // ��ϣ����ʽ
    output              wire   [15:0]                           o_hash_init_val_regs_3             , // ��ϣ����ʽ��ʼֵ
    output              wire                                    o_hash_regs_vld_3                  ,
    output              wire                                    o_port_rxmac_down_regs_3           , // �˿ڽ��շ���MAC�ر�ʹ��
    output              wire                                    o_port_broadcast_drop_regs_3       , // �˿ڹ㲥֡����ʹ��
    output              wire                                    o_port_multicast_drop_regs_3       , // �˿��鲥֡����ʹ��
    output              wire                                    o_port_loopback_drop_regs_3        , // �˿ڻ���֡����ʹ��
    output              wire   [47:0]                           o_port_mac_regs_3                  , // �˿ڵ� MAC ��ַ
    output              wire                                    o_port_mac_vld_regs_3              , // ʹ�ܶ˿� MAC ��ַ��Ч
    output              wire   [7:0]                            o_port_mtu_regs_3                  , // MTU����ֵ
    output              wire   [PORT_NUM-1:0]                   o_port_mirror_frwd_regs_3          , // ����ת���Ĵ���������Ӧ�Ķ˿���1���򱾶˿ڽ��յ����κ�ת������֡������ת��ֵ����1�Ķ˿�
    output              wire   [15:0]                           o_port_flowctrl_cfg_regs_3         , // ������������
    output              wire   [4:0]                            o_port_rx_ultrashortinterval_num_3 , // ֡���
    // ACL �Ĵ�
    output              wire   [PORT_NUM-1:0]                   o_acl_port_sel_3                    , // ѡ��Ҫ���õĶ˿�
    output              wire                                    o_acl_clr_list_regs_3               , // ��ռĴ����б�
    input               wire                                    i_acl_list_rdy_regs_3               , // ���üĴ�����������
    output              wire   [4:0]                            o_acl_item_sel_regs_3               , // ������Ŀѡ��
    //output              wire   [5:0]                            o_acl_item_waddr_regs_3             , // ÿ����Ŀ���֧�ֱȶ� 64 �ֽ�
    //output              wire   [7:0]                            o_acl_item_din_regs_3               , // ��Ҫ�Ƚϵ��ֽ�����
    //output              wire                                    o_acl_item_we_regs_3                , // ����ʹ���ź�
    //output              wire   [15:0]                           o_acl_item_rslt_regs_3              , // ƥ��Ľ��ֵ - [7:0] ���֡����, [15:8] ACLת��ָ���˿�
    //output              wire                                    o_acl_item_complete_regs_3          , // �˿� ACL �����������ʹ���ź�
    output              wire   [95:0]                           o_acl_item_dmac_code_3                ,
    output              wire   [95:0]                           o_acl_item_smac_code_3                ,
    output              wire   [63:0]                           o_acl_item_vlan_code_3                ,
    output              wire   [31:0]                           o_acl_item_ethtype_code_3             ,
    output              wire   [5:0]                            o_acl_item_action_pass_state_3        ,
    output              wire   [15:0]                           o_acl_item_action_cb_streamhandle_3   ,
    output              wire   [5:0]                            o_acl_item_action_flowctrl_3          ,
    output              wire   [15:0]                           o_acl_item_action_txport_3            ,
    // ״̬�Ĵ���
    input              wire   [15:0]                            i_port_diag_state_3                 , // �˿�״̬�Ĵ�����������Ĵ�����˵������ 
    // ��ϼĴ���
    input              wire                                     i_port_rx_ultrashort_frm_3          , // �˿ڽ��ճ���֡(С��64�ֽ�)
    input              wire                                     i_port_rx_overlength_frm_3          , // �˿ڽ��ճ���֡(����MTU�ֽ�)
    input              wire                                     i_port_rx_crcerr_frm_3              , // �˿ڽ���CRC����֡
    input              wire  [15:0]                             i_port_rx_loopback_frm_cnt_3        , // �˿ڽ��ջ���֡������ֵ
    input              wire  [15:0]                             i_port_broadflow_drop_cnt_3         , // �˿ڽ��յ��㲥������������֡������ֵ
    input              wire  [15:0]                             i_port_multiflow_drop_cnt_3         , // �˿ڽ��յ��鲥������������֡������ֵ
    // ����ͳ�ƼĴ���
    input              wire  [15:0]                             i_port_rx_byte_cnt_3                , // �˿�0�����ֽڸ���������ֵ
    input              wire  [15:0]                             i_port_rx_frame_cnt_3               ,  // �˿�0����֡����������ֵ 

    //qbu_rx�Ĵ���  
    input              wire                                     i_rx_busy_3                          , // ����æ�ź�
    input              wire  [15:0]                             i_rx_fragment_cnt_3                  , // ���շ�Ƭ����
    input              wire                                     i_rx_fragment_mismatch_3             , // ��Ƭ��ƥ��
    input              wire  [15:0]                             i_err_rx_crc_cnt_3                   , // CRC�������
    input              wire  [15:0]                             i_err_rx_frame_cnt_3                 , // ֡�������
    input              wire  [15:0]                             i_err_fragment_cnt_3                 , // ��Ƭ�������
    input              wire  [15:0]                             i_rx_frames_cnt_3                    , // ����֡����
    input              wire  [7:0]                              i_frag_next_rx_3                     , // ��һ����Ƭ��
    input              wire  [7:0]                              i_frame_seq_3                        , // ֡���
    output             wire                                     o_reset_3                            ,
`endif
`ifdef MAC4
    output              wire   [15:0]                           o_hash_ploy_regs_4                 , // ��ϣ����ʽ
    output              wire   [15:0]                           o_hash_init_val_regs_4             , // ��ϣ����ʽ��ʼֵ
    output              wire                                    o_hash_regs_vld_4                  ,
    output              wire                                    o_port_rxmac_down_regs_4           , // �˿ڽ��շ���MAC�ر�ʹ��
    output              wire                                    o_port_broadcast_drop_regs_4       , // �˿ڹ㲥֡����ʹ��
    output              wire                                    o_port_multicast_drop_regs_4       , // �˿��鲥֡����ʹ��
    output              wire                                    o_port_loopback_drop_regs_4        , // �˿ڻ���֡����ʹ��
    output              wire   [47:0]                           o_port_mac_regs_4                  , // �˿ڵ� MAC ��ַ
    output              wire                                    o_port_mac_vld_regs_4              , // ʹ�ܶ˿� MAC ��ַ��Ч
    output              wire   [7:0]                            o_port_mtu_regs_4                  , // MTU����ֵ
    output              wire   [PORT_NUM-1:0]                   o_port_mirror_frwd_regs_4          , // ����ת���Ĵ���������Ӧ�Ķ˿���1���򱾶˿ڽ��յ����κ�ת������֡������ת��ֵ����1�Ķ˿�
    output              wire   [15:0]                           o_port_flowctrl_cfg_regs_4         , // ������������
    output              wire   [4:0]                            o_port_rx_ultrashortinterval_num_4 , // ֡���
    // ACL �Ĵ�
    output              wire   [PORT_NUM-1:0]                   o_acl_port_sel_4                    , // ѡ��Ҫ���õĶ˿�
    output              wire                                    o_acl_clr_list_regs_4               , // ��ռĴ����б�
    input               wire                                    i_acl_list_rdy_regs_4               , // ���üĴ�����������
    output              wire   [4:0]                            o_acl_item_sel_regs_4               , // ������Ŀѡ��
    //output              wire   [5:0]                            o_acl_item_waddr_regs_4             , // ÿ����Ŀ���֧�ֱȶ� 64 �ֽ�
    //output              wire   [7:0]                            o_acl_item_din_regs_4               , // ��Ҫ�Ƚϵ��ֽ�����
    //output              wire                                    o_acl_item_we_regs_4                , // ����ʹ���ź�
    //output              wire   [15:0]                           o_acl_item_rslt_regs_4              , // ƥ��Ľ��ֵ - [7:0] ���֡����, [15:8] ACLת��ָ���˿�
    //output              wire                                    o_acl_item_complete_regs_4          , // �˿� ACL �����������ʹ���ź�
    output              wire   [95:0]                           o_acl_item_dmac_code_4                ,
    output              wire   [95:0]                           o_acl_item_smac_code_4                ,
    output              wire   [63:0]                           o_acl_item_vlan_code_4                ,
    output              wire   [31:0]                           o_acl_item_ethtype_code_4             ,
    output              wire   [5:0]                            o_acl_item_action_pass_state_4        ,
    output              wire   [15:0]                           o_acl_item_action_cb_streamhandle_4   ,
    output              wire   [5:0]                            o_acl_item_action_flowctrl_4          ,
    output              wire   [15:0]                           o_acl_item_action_txport_4            ,
    // ״̬�Ĵ���
    input              wire   [15:0]                            i_port_diag_state_4                 , // �˿�״̬�Ĵ�����������Ĵ�����˵������ 
    // ��ϼĴ���
    input              wire                                     i_port_rx_ultrashort_frm_4          , // �˿ڽ��ճ���֡(С��64�ֽ�)
    input              wire                                     i_port_rx_overlength_frm_4          , // �˿ڽ��ճ���֡(����MTU�ֽ�)
    input              wire                                     i_port_rx_crcerr_frm_4              , // �˿ڽ���CRC����֡
    input              wire  [15:0]                             i_port_rx_loopback_frm_cnt_4        , // �˿ڽ��ջ���֡������ֵ
    input              wire  [15:0]                             i_port_broadflow_drop_cnt_4         , // �˿ڽ��յ��㲥������������֡������ֵ
    input              wire  [15:0]                             i_port_multiflow_drop_cnt_4         , // �˿ڽ��յ��鲥������������֡������ֵ
    // ����ͳ�ƼĴ���
    input              wire  [15:0]                             i_port_rx_byte_cnt_4                , // �˿�0�����ֽڸ���������ֵ
    input              wire  [15:0]                             i_port_rx_frame_cnt_4               ,  // �˿�0����֡����������ֵ  

    //qbu_rx�Ĵ���  
    input              wire                                     i_rx_busy_4                          , // ����æ�ź�
    input              wire  [15:0]                             i_rx_fragment_cnt_4                  , // ���շ�Ƭ����
    input              wire                                     i_rx_fragment_mismatch_4             , // ��Ƭ��ƥ��
    input              wire  [15:0]                             i_err_rx_crc_cnt_4                   , // CRC�������
    input              wire  [15:0]                             i_err_rx_frame_cnt_4                 , // ֡�������
    input              wire  [15:0]                             i_err_fragment_cnt_4                 , // ��Ƭ�������
    input              wire  [15:0]                             i_rx_frames_cnt_4                    , // ����֡����
    input              wire  [7:0]                              i_frag_next_rx_4                     , // ��һ����Ƭ��
    input              wire  [7:0]                              i_frame_seq_4                        , // ֡���
    output             wire                                     o_reset_4                            ,
`endif
`ifdef MAC5
    output              wire   [15:0]                           o_hash_ploy_regs_5                 , // ��ϣ����ʽ
    output              wire   [15:0]                           o_hash_init_val_regs_5             , // ��ϣ����ʽ��ʼֵ
    output              wire                                    o_hash_regs_vld_5                  ,
    output              wire                                    o_port_rxmac_down_regs_5           , // �˿ڽ��շ���MAC�ر�ʹ��
    output              wire                                    o_port_broadcast_drop_regs_5       , // �˿ڹ㲥֡����ʹ��
    output              wire                                    o_port_multicast_drop_regs_5       , // �˿��鲥֡����ʹ��
    output              wire                                    o_port_loopback_drop_regs_5        , // �˿ڻ���֡����ʹ��
    output              wire   [47:0]                           o_port_mac_regs_5                  , // �˿ڵ� MAC ��ַ
    output              wire                                    o_port_mac_vld_regs_5              , // ʹ�ܶ˿� MAC ��ַ��Ч
    output              wire   [7:0]                            o_port_mtu_regs_5                  , // MTU����ֵ
    output              wire   [PORT_NUM-1:0]                   o_port_mirror_frwd_regs_5          , // ����ת���Ĵ���������Ӧ�Ķ˿���1���򱾶˿ڽ��յ����κ�ת������֡������ת��ֵ����1�Ķ˿�
    output              wire   [15:0]                           o_port_flowctrl_cfg_regs_5         , // ������������
    output              wire   [4:0]                            o_port_rx_ultrashortinterval_num_5 , // ֡���
    // ACL �Ĵ�
    output              wire   [PORT_NUM-1:0]                   o_acl_port_sel_5                    , // ѡ��Ҫ���õĶ˿�
    output              wire                                    o_acl_clr_list_regs_5               , // ��ռĴ����б�
    input               wire                                    i_acl_list_rdy_regs_5               , // ���üĴ�����������
    output              wire   [4:0]                            o_acl_item_sel_regs_5               , // ������Ŀѡ��
    //output              wire   [5:0]                            o_acl_item_waddr_regs_5             , // ÿ����Ŀ���֧�ֱȶ� 64 �ֽ�
    //output              wire   [7:0]                            o_acl_item_din_regs_5               , // ��Ҫ�Ƚϵ��ֽ�����
    //output              wire                                    o_acl_item_we_regs_5                , // ����ʹ���ź�
    //output              wire   [15:0]                           o_acl_item_rslt_regs_5              , // ƥ��Ľ��ֵ - [7:0] ���֡����, [15:8] ACLת��ָ���˿�
    //output              wire                                    o_acl_item_complete_regs_5          , // �˿� ACL �����������ʹ���ź�
    output              wire   [95:0]                           o_acl_item_dmac_code_5                ,
    output              wire   [95:0]                           o_acl_item_smac_code_5                ,
    output              wire   [63:0]                           o_acl_item_vlan_code_5                ,
    output              wire   [31:0]                           o_acl_item_ethtype_code_5             ,
    output              wire   [5:0]                            o_acl_item_action_pass_state_5        ,
    output              wire   [15:0]                           o_acl_item_action_cb_streamhandle_5   ,
    output              wire   [5:0]                            o_acl_item_action_flowctrl_5          ,
    output              wire   [15:0]                           o_acl_item_action_txport_5            ,
    // ״̬�Ĵ���
    input              wire   [15:0]                            i_port_diag_state_5                 , // �˿�״̬�Ĵ�����������Ĵ�����˵������ 
    // ��ϼĴ���
    input              wire                                     i_port_rx_ultrashort_frm_5          , // �˿ڽ��ճ���֡(С��64�ֽ�)
    input              wire                                     i_port_rx_overlength_frm_5          , // �˿ڽ��ճ���֡(����MTU�ֽ�)
    input              wire                                     i_port_rx_crcerr_frm_5              , // �˿ڽ���CRC����֡
    input              wire  [15:0]                             i_port_rx_loopback_frm_cnt_5        , // �˿ڽ��ջ���֡������ֵ
    input              wire  [15:0]                             i_port_broadflow_drop_cnt_5         , // �˿ڽ��յ��㲥������������֡������ֵ
    input              wire  [15:0]                             i_port_multiflow_drop_cnt_5         , // �˿ڽ��յ��鲥������������֡������ֵ
    // ����ͳ�ƼĴ���
    input              wire  [15:0]                             i_port_rx_byte_cnt_5                , // �˿�0�����ֽڸ���������ֵ
    input              wire  [15:0]                             i_port_rx_frame_cnt_5               ,  // �˿�0����֡����������ֵ  

    //qbu_rx�Ĵ���  
    input              wire                                     i_rx_busy_5                          , // ����æ�ź�
    input              wire  [15:0]                             i_rx_fragment_cnt_5                  , // ���շ�Ƭ����
    input              wire                                     i_rx_fragment_mismatch_5             , // ��Ƭ��ƥ��
    input              wire  [15:0]                             i_err_rx_crc_cnt_5                   , // CRC�������
    input              wire  [15:0]                             i_err_rx_frame_cnt_5                 , // ֡�������
    input              wire  [15:0]                             i_err_fragment_cnt_5                 , // ��Ƭ�������
    input              wire  [15:0]                             i_rx_frames_cnt_5                    , // ����֡����
    input              wire  [7:0]                              i_frag_next_rx_5                     , // ��һ����Ƭ��
    input              wire  [7:0]                              i_frame_seq_5                        , // ֡���
    output             wire                                     o_reset_5                            ,
`endif
`ifdef MAC6
    output              wire   [15:0]                           o_hash_ploy_regs_6                 , // ��ϣ����ʽ
    output              wire   [15:0]                           o_hash_init_val_regs_6             , // ��ϣ����ʽ��ʼֵ
    output              wire                                    o_hash_regs_vld_6                  ,
    output              wire                                    o_port_rxmac_down_regs_6           , // �˿ڽ��շ���MAC�ر�ʹ��
    output              wire                                    o_port_broadcast_drop_regs_6       , // �˿ڹ㲥֡����ʹ��
    output              wire                                    o_port_multicast_drop_regs_6       , // �˿��鲥֡����ʹ��
    output              wire                                    o_port_loopback_drop_regs_6        , // �˿ڻ���֡����ʹ��
    output              wire   [47:0]                           o_port_mac_regs_6                  , // �˿ڵ� MAC ��ַ
    output              wire                                    o_port_mac_vld_regs_6              , // ʹ�ܶ˿� MAC ��ַ��Ч
    output              wire   [7:0]                            o_port_mtu_regs_6                  , // MTU����ֵ
    output              wire   [PORT_NUM-1:0]                   o_port_mirror_frwd_regs_6          , // ����ת���Ĵ���������Ӧ�Ķ˿���1���򱾶˿ڽ��յ����κ�ת������֡������ת��ֵ����1�Ķ˿�
    output              wire   [15:0]                           o_port_flowctrl_cfg_regs_6         , // ������������
    output              wire   [4:0]                            o_port_rx_ultrashortinterval_num_6 , // ֡���
    // ACL �Ĵ�
    output              wire   [PORT_NUM-1:0]                   o_acl_port_sel_6                    , // ѡ��Ҫ���õĶ˿�
    output              wire                                    o_acl_clr_list_regs_6               , // ��ռĴ����б�
    input               wire                                    i_acl_list_rdy_regs_6               , // ���üĴ�����������
    output              wire   [4:0]                            o_acl_item_sel_regs_6               , // ������Ŀѡ��
    //output              wire   [5:0]                            o_acl_item_waddr_regs_6             , // ÿ����Ŀ���֧�ֱȶ� 64 �ֽ�
    //output              wire   [7:0]                            o_acl_item_din_regs_6               , // ��Ҫ�Ƚϵ��ֽ�����
    //output              wire                                    o_acl_item_we_regs_6                , // ����ʹ���ź�
    //output              wire   [15:0]                           o_acl_item_rslt_regs_6              , // ƥ��Ľ��ֵ - [7:0] ���֡����, [15:8] ACLת��ָ���˿�
    //output              wire                                    o_acl_item_complete_regs_6          , // �˿� ACL �����������ʹ���ź�
    output              wire   [95:0]                           o_acl_item_dmac_code_6                ,
    output              wire   [95:0]                           o_acl_item_smac_code_6                ,
    output              wire   [63:0]                           o_acl_item_vlan_code_6                ,
    output              wire   [31:0]                           o_acl_item_ethtype_code_6             ,
    output              wire   [5:0]                            o_acl_item_action_pass_state_6        ,
    output              wire   [15:0]                           o_acl_item_action_cb_streamhandle_6   ,
    output              wire   [5:0]                            o_acl_item_action_flowctrl_6          ,
    output              wire   [15:0]                           o_acl_item_action_txport_6            ,
    // ״̬�Ĵ���
    input              wire   [15:0]                            i_port_diag_state_6                 , // �˿�״̬�Ĵ�����������Ĵ�����˵������ 
    // ��ϼĴ���
    input              wire                                     i_port_rx_ultrashort_frm_6          , // �˿ڽ��ճ���֡(С��64�ֽ�)
    input              wire                                     i_port_rx_overlength_frm_6          , // �˿ڽ��ճ���֡(����MTU�ֽ�)
    input              wire                                     i_port_rx_crcerr_frm_6              , // �˿ڽ���CRC����֡
    input              wire  [15:0]                             i_port_rx_loopback_frm_cnt_6        , // �˿ڽ��ջ���֡������?
    input              wire  [15:0]                             i_port_broadflow_drop_cnt_6         , // �˿ڽ��յ��㲥������������֡������ֵ
    input              wire  [15:0]                             i_port_multiflow_drop_cnt_6         , // �˿ڽ��յ��鲥������������֡������?
    // ����ͳ�ƼĴ���
    input              wire  [15:0]                             i_port_rx_byte_cnt_6                , // �˿�0�����ֽڸ���������ֵ
    input              wire  [15:0]                             i_port_rx_frame_cnt_6               ,  // �˿�0����֡����������ֵ  

    //qbu_rx�Ĵ���  
    input              wire                                     i_rx_busy_6                          , // ����æ�ź�
    input              wire  [15:0]                             i_rx_fragment_cnt_6                  , // ���շ�Ƭ����
    input              wire                                     i_rx_fragment_mismatch_6             , // ��Ƭ��ƥ��
    input              wire  [15:0]                             i_err_rx_crc_cnt_6                   , // CRC�������
    input              wire  [15:0]                             i_err_rx_frame_cnt_6                 , // ֡�������
    input              wire  [15:0]                             i_err_fragment_cnt_6                 , // ��Ƭ�������
    input              wire  [15:0]                             i_rx_frames_cnt_6                    , // ����֡����
    input              wire  [7:0]                              i_frag_next_rx_6                     , // ��һ����Ƭ��
    input              wire  [7:0]                              i_frame_seq_6                        , // ֡���
    output             wire                                     o_reset_6                            ,
`endif
`ifdef MAC7
    output              wire   [15:0]                           o_hash_ploy_regs_7                , // ��ϣ����ʽ
    output              wire   [15:0]                           o_hash_init_val_regs_7            , // ��ϣ����ʽ��ʼֵ
    output              wire                                    o_hash_regs_vld_7                 ,
    output              wire                                    o_port_rxmac_down_regs_7          , // �˿ڽ��շ���MAC�ر�ʹ��
    output              wire                                    o_port_broadcast_drop_regs_7      , // �˿ڹ㲥֡����ʹ��
    output              wire                                    o_port_multicast_drop_regs_7      , // �˿��鲥֡����ʹ��
    output              wire                                    o_port_loopback_drop_regs_7       , // �˿ڻ���֡����ʹ��
    output              wire   [47:0]                           o_port_mac_regs_7                 , // �˿ڵ� MAC ��ַ
    output              wire                                    o_port_mac_vld_regs_7             , // ʹ�ܶ˿� MAC ��ַ��Ч
    output              wire   [7:0]                            o_port_mtu_regs_7                 , // MTU����ֵ
    output              wire   [PORT_NUM-1:0]                   o_port_mirror_frwd_regs_7         , // ����ת���Ĵ���������Ӧ�Ķ˿���1���򱾶˿ڽ��յ����κ�ת������֡������ת��ֵ����1�Ķ˿�
    output              wire   [15:0]                           o_port_flowctrl_cfg_regs_7        , // ������������
    output              wire   [4:0]                            o_port_rx_ultrashortinterval_num_7, // ֡���
    // ACL �Ĵ�
    output              wire   [PORT_NUM-1:0]                   o_acl_port_sel_7                   , // ѡ��Ҫ���õĶ˿�
    output              wire                                    o_acl_clr_list_regs_7              , // ��ռĴ����б�
    input               wire                                    i_acl_list_rdy_regs_7              , // ���üĴ�����������
    output              wire   [4:0]                            o_acl_item_sel_regs_7              , // ������Ŀѡ��
    //output              wire   [5:0]                            o_acl_item_waddr_regs_7            , // ÿ����Ŀ���֧�ֱȶ� 64 �ֽ�
    //output              wire   [7:0]                            o_acl_item_din_regs_7              , // ��Ҫ�Ƚϵ��ֽ�����
    //output              wire                                    o_acl_item_we_regs_7               , // ����ʹ���ź�
    //output              wire   [15:0]                           o_acl_item_rslt_regs_7             , // ƥ��Ľ��ֵ - [7:0] ���֡����, [15:8] ACLת��ָ���˿�
    //output              wire                                    o_acl_item_complete_regs_7         , // �˿� ACL �����������ʹ���ź�
    output              wire   [95:0]                           o_acl_item_dmac_code_7                ,
    output              wire   [95:0]                           o_acl_item_smac_code_7                ,
    output              wire   [63:0]                           o_acl_item_vlan_code_7                ,
    output              wire   [31:0]                           o_acl_item_ethtype_code_7             ,
    output              wire   [5:0]                            o_acl_item_action_pass_state_7        ,
    output              wire   [15:0]                           o_acl_item_action_cb_streamhandle_7   ,
    output              wire   [5:0]                            o_acl_item_action_flowctrl_7          ,
    output              wire   [15:0]                           o_acl_item_action_txport_7            ,
    // ״̬�Ĵ���
    input              wire   [15:0]                            i_port_diag_state_7                , // �˿�״̬�Ĵ�����������Ĵ�����˵������ 
    // ��ϼĴ���
    input              wire                                     i_port_rx_ultrashort_frm_7         , // �˿ڽ��ճ���֡(С��64�ֽ�)
    input              wire                                     i_port_rx_overlength_frm_7         , // �˿ڽ��ճ���֡(����MTU�ֽ�)
    input              wire                                     i_port_rx_crcerr_frm_7             , // �˿ڽ���CRC����֡
    input              wire  [15:0]                             i_port_rx_loopback_frm_cnt_7       , // �˿ڽ��ջ���֡������ֵ
    input              wire  [15:0]                             i_port_broadflow_drop_cnt_7        , // �˿ڽ��յ��㲥������������֡������ֵ
    input              wire  [15:0]                             i_port_multiflow_drop_cnt_7        , // �˿ڽ��յ��鲥������������֡������?
    // ����ͳ�ƼĴ���
    input              wire  [15:0]                             i_port_rx_byte_cnt_7               , // �˿�0�����ֽڸ���������ֵ
    input              wire  [15:0]                             i_port_rx_frame_cnt_7              , // �˿�0����֡����������ֵ  

    //qbu_rx�Ĵ���  
    input              wire                                     i_rx_busy_7                          , // ����æ�ź�
    input              wire  [15:0]                             i_rx_fragment_cnt_7                  , // ���շ�Ƭ����
    input              wire                                     i_rx_fragment_mismatch_7             , // ��Ƭ��ƥ��
    input              wire  [15:0]                             i_err_rx_crc_cnt_7                   , // CRC�������
    input              wire  [15:0]                             i_err_rx_frame_cnt_7                 , // ֡�������
    input              wire  [15:0]                             i_err_fragment_cnt_7                 , // ��Ƭ�������
    input              wire  [15:0]                             i_rx_frames_cnt_7                    , // ����֡����
    input              wire  [7:0]                              i_frag_next_rx_7                     , // ��һ����Ƭ��
    input              wire  [7:0]                              i_frame_seq_7                        , // ֡���
    output             wire                                     o_reset_7                            ,
`endif
    /*---------------------------------------- �Ĵ������ýӿ� -------------------------------------------*/
    // �Ĵ��������ź�                     
    input              wire                                     i_refresh_list_pulse                , // ˢ�¼Ĵ����б�״̬�Ĵ����Ϳ��ƼĴ�����
    input              wire                                     i_switch_err_cnt_clr                , // ˢ�´��������
    input              wire                                     i_switch_err_cnt_stat               , // ˢ�´���״̬�Ĵ���
    // �Ĵ���д���ƽӿ�     
    input              wire                                     i_switch_reg_bus_we                 , // �Ĵ���дʹ��
    input              wire   [REG_ADDR_BUS_WIDTH-1:0]          i_switch_reg_bus_we_addr            , // �Ĵ���д��ַ
    input              wire   [REG_DATA_BUS_WIDTH-1:0]          i_switch_reg_bus_we_din             , // �Ĵ���д����
    input              wire                                     i_switch_reg_bus_we_din_v           , // �Ĵ���д����ʹ��
    // �Ĵ��������ƽӿ�     
    input              wire                                     i_switch_reg_bus_rd                 , // �Ĵ�����ʹ��
    input              wire   [REG_ADDR_BUS_WIDTH-1:0]          i_switch_reg_bus_rd_addr            , // �Ĵ�������ַ
    output             wire   [REG_DATA_BUS_WIDTH-1:0]          o_switch_reg_bus_rd_dout            , // �����Ĵ�������
    output             wire                                     o_switch_reg_bus_rd_dout_v           // ��������Чʹ��
);

/*---------------------------------------- RXMAC�Ĵ�����ַ���� -------------------------------------------*/
localparam  REG_HASH_PLOY                   		=   8'h00                   ;
localparam  REG_HASH_INIT_VAL               		=   8'h01                   ;
localparam  REG_PORT_RXMAC_DOWN            	 		=   8'h02                   ;
localparam  REG_PORT_ACL_ENABLE             		=	8'h03					;
localparam  REG_PORT_BROADCAST_DROP         		=   8'h04					;
localparam  REG_PORT_MULTICAST_DROP                 =   8'h05					;
localparam  REG_PORT_LOOKBACK_DROP                  =   8'h06					;
localparam  REG_PORT_FORCE_RECAL_CRC                =   8'h07					;
localparam  REG_PORT_FLOODFRM_DROP                  =   8'h08					;
localparam  REG_PORT_MULTIFLOOD_DROP                =   8'h09					;
localparam  REG_CFG_RXMAC_PORT_SEL                  =   8'h10					;
localparam  REG_PORTMTU                             =   8'h11					;
localparam  REG_PORTMAC0                            =   8'h12					;
localparam  REG_PORTMAC1                            =   8'h13					;
localparam  REG_PORTMAC2                            =   8'h14					;
localparam  REG_PORTMAC_VALID                       =   8'h15					;
localparam  REG_PORT_MIRROR_FRWD                    =   8'h16					;
localparam  REG_PORT_FLOWCTRL_CFG                   =   8'h17					;
localparam  REG_CFG_ACL_PORT_SEL                    =   8'h20					;
localparam  REG_CFG_ACL_CLR_LIST                    =   8'h21					;
localparam  REG_CFG_ACL_LIST_RDY                    =   8'h22					;
localparam  REG_CFG_ACL_ITEM_SEL                    =   8'h23					;
localparam  REG_CFG_ACL_ITEM_DMAC_CODE_1            =   8'h24					;
localparam  REG_CFG_ACL_ITEM_DMAC_CODE_2            =   8'h25					;
localparam  REG_CFG_ACL_ITEM_DMAC_CODE_3            =   8'h26					;
localparam  REG_CFG_ACL_ITEM_DMAC_CODE_4            =   8'h27					;
localparam  REG_CFG_ACL_ITEM_DMAC_CODE_5            =   8'h28					;
localparam  REG_CFG_ACL_ITEM_DMAC_CODE_6            =   8'h29					;
localparam  REG_CFG_ACL_ITEM_SMAC_CODE_1            =   8'h2A					;
localparam  REG_CFG_ACL_ITEM_SMAC_CODE_2            =   8'h2B					;
localparam  REG_CFG_ACL_ITEM_SMAC_CODE_3            =   8'h2C					;
localparam  REG_CFG_ACL_ITEM_SMAC_CODE_4            =   8'h2D					;
localparam  REG_CFG_ACL_ITEM_SMAC_CODE_5            =   8'h2E					;
localparam  REG_CFG_ACL_ITEM_SMAC_CODE_6            =   8'h2F					;
localparam  REG_CFG_ACL_ITEM_VLAN_CODE_1            =   8'h30					;
localparam  REG_CFG_ACL_ITEM_VLAN_CODE_2            =   8'h31					;
localparam  REG_CFG_ACL_ITEM_VLAN_CODE_3            =   8'h32					;
localparam  REG_CFG_ACL_ITEM_VLAN_CODE_4            =   8'h33					;
localparam  REG_CFG_ACL_ITEM_ETHTYPE_CODE_1         =   8'h34					;
localparam  REG_CFG_ACL_ITEM_ETHTYPE_CODE_2         =   8'h35					;
localparam  REG_CFG_ACL_ITEM_ACTION_PASS_STATE      =   8'h36					;
localparam  REG_CFG_ACL_ITEM_ACTION_CB_STREAMHANDLE =   8'h37					;
localparam  REG_CFG_ACL_ITEM_ACTION_FLOWCTRL		=   8'h38					;
localparam  REG_CFG_ACL_ITEM_ACTION_TXPORT			=   8'h39					;																
localparam  REG_PORT_RX_BYTE_CNT_0					=   8'h50					;
localparam  REG_PORT_RX_FRAME_CNT_0                 =   8'h51					;
localparam  REG_PORT_DIAG_STATE_0                   =   8'h52					;
localparam  REG_PORT_RX_ULTRASHORT_FRM_CNT_0        =   8'h53					;
localparam  REG_PORT_RX_OVERLENGTH_FRM_CNT_0        =   8'h54					;
localparam  REG_PORT_RX_CRCERR_FRM_CNT_0            =   8'h55					;
localparam  REG_PORT_RX_LOOKBACK_FRM_CNT_0          =   8'h56					;
localparam  REG_PORT_RX_ERROR_DROP_CNT_0            =   8'h57					;
localparam  REG_PORT_BROADFLOW_DROP_CNT_0           =   8'h58					;
localparam  REG_PORT_MULTIFLOW_DROP_CNT_0           =   8'h59					;
localparam  REG_PORT_FLOODFLOW_DROP_CNT_0           =   8'h5A					;
localparam  REG_PORT_RX_OVERPREMB_FRM_CNT_0         =   8'h5B					;
localparam  REG_PORT_RX_ULTRASHORTPREMB_NUM_0       =   8'h5C					;
localparam  REG_PORT_RX_ULTRASHORTINTERVAL_NUM_0    =   8'h5D					;
localparam  REG_PORT_RX_ERRORPREMB_FRM_CNT_0        =   8'h5E					;
localparam  REG_PORT_RX_BYTE_CNT_1					=   8'h60					;
localparam  REG_PORT_RX_FRAME_CNT_1                 =   8'h61					;
localparam  REG_PORT_DIAG_STATE_1                   =   8'h62					;
localparam  REG_PORT_RX_ULTRASHORT_FRM_CNT_1        =   8'h63					;
localparam  REG_PORT_RX_OVERLENGTH_FRM_CNT_1        =   8'h64					;
localparam  REG_PORT_RX_CRCERR_FRM_CNT_1            =   8'h65					;
localparam  REG_PORT_RX_LOOKBACK_FRM_CNT_1          =   8'h66					;
localparam  REG_PORT_RX_ERROR_DROP_CNT_1            =   8'h67					;
localparam  REG_PORT_BROADFLOW_DROP_CNT_1           =   8'h68					;
localparam  REG_PORT_MULTIFLOW_DROP_CNT_1           =   8'h69					;
localparam  REG_PORT_FLOODFLOW_DROP_CNT_1           =   8'h6A					;
localparam  REG_PORT_RX_OVERPREMB_FRM_CNT_1         =   8'h6B					;
localparam  REG_PORT_RX_ULTRASHORTPREMB_NUM_1       =   8'h6C					;
localparam  REG_PORT_RX_ULTRASHORTINTERVAL_NUM_1    =   8'h6D					;
localparam  REG_PORT_RX_ERRORPREMB_FRM_CNT_1        =   8'h6E					;
localparam  REG_PORT_RX_BYTE_CNT_2					=   8'h70					;
localparam  REG_PORT_RX_FRAME_CNT_2                 =   8'h71					;
localparam  REG_PORT_DIAG_STATE_2                   =   8'h72					;
localparam  REG_PORT_RX_ULTRASHORT_FRM_CNT_2        =   8'h73					;
localparam  REG_PORT_RX_OVERLENGTH_FRM_CNT_2        =   8'h74					;
localparam  REG_PORT_RX_CRCERR_FRM_CNT_2            =   8'h75					;
localparam  REG_PORT_RX_LOOKBACK_FRM_CNT_2          =   8'h76					;
localparam  REG_PORT_RX_ERROR_DROP_CNT_2            =   8'h77					;
localparam  REG_PORT_BROADFLOW_DROP_CNT_2           =   8'h78					;
localparam  REG_PORT_MULTIFLOW_DROP_CNT_2           =   8'h79					;
localparam  REG_PORT_FLOODFLOW_DROP_CNT_2           =   8'h7A					;
localparam  REG_PORT_RX_OVERPREMB_FRM_CNT_2         =   8'h7B					;
localparam  REG_PORT_RX_ULTRASHORTPREMB_NUM_2       =   8'h7C					;
localparam  REG_PORT_RX_ULTRASHORTINTERVAL_NUM_2    =   8'h7D					;
localparam  REG_PORT_RX_ERRORPREMB_FRM_CNT_2        =   8'h7E					;
localparam  REG_PORT_RX_BYTE_CNT_3					=   8'h80					;
localparam  REG_PORT_RX_FRAME_CNT_3                 =   8'h81					;
localparam  REG_PORT_DIAG_STATE_3                   =   8'h82					;
localparam  REG_PORT_RX_ULTRASHORT_FRM_CNT_3        =   8'h83					;
localparam  REG_PORT_RX_OVERLENGTH_FRM_CNT_3        =   8'h84					;
localparam  REG_PORT_RX_CRCERR_FRM_CNT_3            =   8'h85					;
localparam  REG_PORT_RX_LOOKBACK_FRM_CNT_3          =   8'h86					;
localparam  REG_PORT_RX_ERROR_DROP_CNT_3            =   8'h87					;
localparam  REG_PORT_BROADFLOW_DROP_CNT_3           =   8'h88					;
localparam  REG_PORT_MULTIFLOW_DROP_CNT_3           =   8'h89					;
localparam  REG_PORT_FLOODFLOW_DROP_CNT_3           =   8'h8A					;
localparam  REG_PORT_RX_OVERPREMB_FRM_CNT_3         =   8'h8B					;
localparam  REG_PORT_RX_ULTRASHORTPREMB_NUM_3       =   8'h8C					;
localparam  REG_PORT_RX_ULTRASHORTINTERVAL_NUM_3    =   8'h8D					;
localparam  REG_PORT_RX_ERRORPREMB_FRM_CNT_3        =   8'h8E					;
localparam  REG_PORT_RX_BYTE_CNT_4					=   8'h90					;
localparam  REG_PORT_RX_FRAME_CNT_4                 =   8'h91					;
localparam  REG_PORT_DIAG_STATE_4                   =   8'h92					;
localparam  REG_PORT_RX_ULTRASHORT_FRM_CNT_4        =   8'h93					;
localparam  REG_PORT_RX_OVERLENGTH_FRM_CNT_4        =   8'h94					;
localparam  REG_PORT_RX_CRCERR_FRM_CNT_4            =   8'h95					;
localparam  REG_PORT_RX_LOOKBACK_FRM_CNT_4          =   8'h96					;
localparam  REG_PORT_RX_ERROR_DROP_CNT_4            =   8'h97					;
localparam  REG_PORT_BROADFLOW_DROP_CNT_4           =   8'h98					;
localparam  REG_PORT_MULTIFLOW_DROP_CNT_4           =   8'h99					;
localparam  REG_PORT_FLOODFLOW_DROP_CNT_4           =   8'h9A					;
localparam  REG_PORT_RX_OVERPREMB_FRM_CNT_4         =   8'h9B					;
localparam  REG_PORT_RX_ULTRASHORTPREMB_NUM_4       =   8'h9C					;
localparam  REG_PORT_RX_ULTRASHORTINTERVAL_NUM_4    =   8'h9D					;
localparam  REG_PORT_RX_ERRORPREMB_FRM_CNT_4        =   8'h9E					;    
localparam  REG_PORT_RX_BYTE_CNT_5					=   8'hA0					;
localparam  REG_PORT_RX_FRAME_CNT_5                 =   8'hA1					;
localparam  REG_PORT_DIAG_STATE_5                   =   8'hA2					;
localparam  REG_PORT_RX_ULTRASHORT_FRM_CNT_5        =   8'hA3					;
localparam  REG_PORT_RX_OVERLENGTH_FRM_CNT_5        =   8'hA4					;
localparam  REG_PORT_RX_CRCERR_FRM_CNT_5            =   8'hA5					;
localparam  REG_PORT_RX_LOOKBACK_FRM_CNT_5          =   8'hA6					;
localparam  REG_PORT_RX_ERROR_DROP_CNT_5            =   8'hA7					;
localparam  REG_PORT_BROADFLOW_DROP_CNT_5           =   8'hA8					;
localparam  REG_PORT_MULTIFLOW_DROP_CNT_5           =   8'hA9					;
localparam  REG_PORT_FLOODFLOW_DROP_CNT_5           =   8'hAA					;
localparam  REG_PORT_RX_OVERPREMB_FRM_CNT_5         =   8'hAB					;
localparam  REG_PORT_RX_ULTRASHORTPREMB_NUM_5       =   8'hAC					;
localparam  REG_PORT_RX_ULTRASHORTINTERVAL_NUM_5    =   8'hAD					;
localparam  REG_PORT_RX_ERRORPREMB_FRM_CNT_5        =   8'hAE					;
localparam  REG_PORT_RX_BYTE_CNT_6					=   8'hB0					;
localparam  REG_PORT_RX_FRAME_CNT_6                 =   8'hB1					;
localparam  REG_PORT_DIAG_STATE_6                   =   8'hB2					;
localparam  REG_PORT_RX_ULTRASHORT_FRM_CNT_6        =   8'hB3					;
localparam  REG_PORT_RX_OVERLENGTH_FRM_CNT_6        =   8'hB4					;
localparam  REG_PORT_RX_CRCERR_FRM_CNT_6            =   8'hB5					;
localparam  REG_PORT_RX_LOOKBACK_FRM_CNT_6          =   8'hB6					;
localparam  REG_PORT_RX_ERROR_DROP_CNT_6            =   8'hB7					;
localparam  REG_PORT_BROADFLOW_DROP_CNT_6           =   8'hB8					;
localparam  REG_PORT_MULTIFLOW_DROP_CNT_6           =   8'hB9					;
localparam  REG_PORT_FLOODFLOW_DROP_CNT_6           =   8'hBA					;
localparam  REG_PORT_RX_OVERPREMB_FRM_CNT_6         =   8'hBB					;
localparam  REG_PORT_RX_ULTRASHORTPREMB_NUM_6       =   8'hBC					;
localparam  REG_PORT_RX_ULTRASHORTINTERVAL_NUM_6    =   8'hBD					;
localparam  REG_PORT_RX_ERRORPREMB_FRM_CNT_6        =   8'hBE					;
localparam  REG_PORT_RX_BYTE_CNT_7					=   8'hC0					;
localparam  REG_PORT_RX_FRAME_CNT_7                 =   8'hC1					;
localparam  REG_PORT_DIAG_STATE_7                   =   8'hC2					;
localparam  REG_PORT_RX_ULTRASHORT_FRM_CNT_7        =   8'hC3					;
localparam  REG_PORT_RX_OVERLENGTH_FRM_CNT_7        =   8'hC4					;
localparam  REG_PORT_RX_CRCERR_FRM_CNT_7            =   8'hC5					;
localparam  REG_PORT_RX_LOOKBACK_FRM_CNT_7          =   8'hC6					;
localparam  REG_PORT_RX_ERROR_DROP_CNT_7            =   8'hC7					;
localparam  REG_PORT_BROADFLOW_DROP_CNT_7           =   8'hC8					;
localparam  REG_PORT_MULTIFLOW_DROP_CNT_7           =   8'hC9					;
localparam  REG_PORT_FLOODFLOW_DROP_CNT_7           =   8'hCA					;
localparam  REG_PORT_RX_OVERPREMB_FRM_CNT_7         =   8'hCB					;
localparam  REG_PORT_RX_ULTRASHORTPREMB_NUM_7       =   8'hCC					;
localparam  REG_PORT_RX_ULTRASHORTINTERVAL_NUM_7    =   8'hCD					;
localparam  REG_PORT_RX_ERRORPREMB_FRM_CNT_7        =   8'hCE					;
/*---------------------------------------- QBU_RX�Ĵ�����ַ���� -------------------------------------------*/
//�˿�1
localparam  REG_QBU_RESET_0                         =   9'hD0                   ;
localparam  REG_RX_FRAGMENT_CNT_0                   =   9'hD1                   ;
localparam  REG_RX_FRAGMENT_MISMATCH_0              =   9'hD2                   ;
localparam  REG_ERR_RX_CRC_CNT_0                    =   9'hD3                   ;
localparam  REG_ERR_RX_FRAME_CNT_0                  =   9'hD4                   ;
localparam  REG_ERR_FRAGMENT_CNT_0                  =   9'hD5                   ;
localparam  REG_ERR_VERIFI_CNT_0                    =   9'hD6                   ;
localparam  REG_RX_FRAMES_CNT_0                     =   9'hD7                   ;
localparam  REG_FRAG_NEXT_RX_0                      =   9'hD8                   ;
localparam  REG_FRAME_SEQ_0                         =   9'hD9                   ;
//�˿�2
localparam  REG_QBU_RESET_1                         =   9'hDA                   ;
localparam  REG_RX_FRAGMENT_CNT_1                   =   9'hDB                   ;
localparam  REG_RX_FRAGMENT_MISMATCH_1              =   9'hDC                   ;
localparam  REG_ERR_RX_CRC_CNT_1                    =   9'hDD                   ;
localparam  REG_ERR_RX_FRAME_CNT_1                  =   9'hDE                   ;
localparam  REG_ERR_FRAGMENT_CNT_1                  =   9'hDF                   ;
localparam  REG_ERR_VERIFI_CNT_1                    =   9'hE0                   ;
localparam  REG_RX_FRAMES_CNT_1                     =   9'hE1                   ;
localparam  REG_FRAG_NEXT_RX_1                      =   9'hE2                   ;
localparam  REG_FRAME_SEQ_1                         =   9'hE3                   ;
//�˿�3
localparam  REG_QBU_RESET_2                         =   9'hE4                   ;
localparam  REG_RX_FRAGMENT_CNT_2                   =   9'hE5                   ;
localparam  REG_RX_FRAGMENT_MISMATCH_2              =   9'hE6                   ;
localparam  REG_ERR_RX_CRC_CNT_2                    =   9'hE7                   ;
localparam  REG_ERR_RX_FRAME_CNT_2                  =   9'hE8                   ;
localparam  REG_ERR_FRAGMENT_CNT_2                  =   9'hE9                   ;
localparam  REG_ERR_VERIFI_CNT_2                    =   9'hEA                   ;
localparam  REG_RX_FRAMES_CNT_2                     =   9'hEB                   ;
localparam  REG_FRAG_NEXT_RX_2                      =   9'hEC                   ;
localparam  REG_FRAME_SEQ_2                         =   9'hED                   ;
//�˿�4
localparam  REG_QBU_RESET_3                         =   9'hEE                   ;
localparam  REG_RX_FRAGMENT_CNT_3                   =   9'hEF                   ;
localparam  REG_RX_FRAGMENT_MISMATCH_3              =   9'hF0                   ;
localparam  REG_ERR_RX_CRC_CNT_3                    =   9'hF1                   ;
localparam  REG_ERR_RX_FRAME_CNT_3                  =   9'hF2                   ;
localparam  REG_ERR_FRAGMENT_CNT_3                  =   9'hF3                   ;
localparam  REG_ERR_VERIFI_CNT_3                    =   9'hF4                   ;
localparam  REG_RX_FRAMES_CNT_3                     =   9'hF5                   ;
localparam  REG_FRAG_NEXT_RX_3                      =   9'hF6                   ;
localparam  REG_FRAME_SEQ_3                         =   9'hF7                   ;
//�˿�5
localparam  REG_QBU_RESET_4                         =   9'hF8                   ;
localparam  REG_RX_FRAGMENT_CNT_4                   =   9'hF9                   ;
localparam  REG_RX_FRAGMENT_MISMATCH_4              =   9'hFA                   ;
localparam  REG_ERR_RX_CRC_CNT_4                    =   9'hFB                   ;
localparam  REG_ERR_RX_FRAME_CNT_4                  =   9'hFC                   ;
localparam  REG_ERR_FRAGMENT_CNT_4                  =   9'hFD                   ;
localparam  REG_ERR_VERIFI_CNT_4                    =   9'hFE                   ;
localparam  REG_RX_FRAMES_CNT_4                     =   9'hFF                   ;
localparam  REG_FRAG_NEXT_RX_4                      =   9'h100                  ;
localparam  REG_FRAME_SEQ_4                         =   9'h101                  ;
//�˿�6
localparam  REG_QBU_RESET_5                         =   9'h102                  ;
localparam  REG_RX_FRAGMENT_CNT_5                   =   9'h103                  ;
localparam  REG_RX_FRAGMENT_MISMATCH_5              =   9'h104                  ;
localparam  REG_ERR_RX_CRC_CNT_5                    =   9'h105                  ;
localparam  REG_ERR_RX_FRAME_CNT_5                  =   9'h106                  ;
localparam  REG_ERR_FRAGMENT_CNT_5                  =   9'h107                  ;
localparam  REG_ERR_VERIFI_CNT_5                    =   9'h108                  ;
localparam  REG_RX_FRAMES_CNT_5                     =   9'h109                  ;
localparam  REG_FRAG_NEXT_RX_5                      =   9'h10A                  ;
localparam  REG_FRAME_SEQ_5                         =   9'h10B                  ;
//�˿�7
localparam  REG_QBU_RESET_6                         =   9'h10C                  ;
localparam  REG_RX_FRAGMENT_CNT_6                   =   9'h10D                  ;
localparam  REG_RX_FRAGMENT_MISMATCH_6              =   9'h10E                  ;
localparam  REG_ERR_RX_CRC_CNT_6                    =   9'h10F                  ;
localparam  REG_ERR_RX_FRAME_CNT_6                  =   9'h110                  ;
localparam  REG_ERR_FRAGMENT_CNT_6                  =   9'h111                  ;
localparam  REG_ERR_VERIFI_CNT_6                    =   9'h112                  ;
localparam  REG_RX_FRAMES_CNT_6                     =   9'h113                  ;
localparam  REG_FRAG_NEXT_RX_6                      =   9'h114                  ;
localparam  REG_FRAME_SEQ_6                         =   9'h115                  ;
//�˿�8
localparam  REG_QBU_RESET_7                         =   9'h116                  ;
localparam  REG_RX_FRAGMENT_CNT_7                   =   9'h117                  ;
localparam  REG_RX_FRAGMENT_MISMATCH_7              =   9'h118                  ;
localparam  REG_ERR_RX_CRC_CNT_7                    =   9'h119                  ;
localparam  REG_ERR_RX_FRAME_CNT_7                  =   9'h11A                  ;
localparam  REG_ERR_FRAGMENT_CNT_7                  =   9'h11B                  ;
localparam  REG_ERR_VERIFI_CNT_7                    =   9'h11C                  ;
localparam  REG_RX_FRAMES_CNT_7                     =   9'h11D                  ;
localparam  REG_FRAG_NEXT_RX_7                      =   9'h11E                  ;
localparam  REG_FRAME_SEQ_7                         =   9'h11F                  ;

/*------------------------------------------- �ڲ��źŶ��� -----------------------------------------------*/
// �Ĵ���ˢ�¿����ź�  
reg                                         r_refresh_list_pulse                ; // ˢ�¼Ĵ����б�״̬�Ĵ����Ϳ��ƼĴ�����
reg                                         r_switch_err_cnt_clr                ; // ˢ�´��������
reg                                         r_switch_err_cnt_stat               ; // ˢ�´���״̬�Ĵ���
/*------------------------------------------- �Ĵ����źŶ��� ------------------------------------------*/
// �Ĵ���д�����ź�  
reg                                         r_reg_bus_we                        ;
reg             [REG_ADDR_BUS_WIDTH-1:0]    r_reg_bus_addr                      ;
reg             [REG_DATA_BUS_WIDTH-1:0]    r_reg_bus_data                      ;
reg                                         r_reg_bus_data_vld                  ;
// �Ĵ����������ź�
reg                                         r_reg_bus_re                        ;
reg             [REG_ADDR_BUS_WIDTH-1:0]    r_reg_bus_raddr                     ;
reg             [REG_DATA_BUS_WIDTH-1:0]    r_reg_bus_rdata                     ;
reg                                         r_reg_bus_rdata_vld                 ;
/*========================================  RXMAC�Ĵ�����д�����źŹ��� ========================================*/
// ͨ�üĴ���
reg   [15:0]                           r_hash_ploy_regs                  ;// ��ϣ����ʽ
reg   [15:0]                           r_hash_init_val_regs              ;// ��ϣ����ʽ��ʼֵ
reg                                    r_hash_regs_vld                   ;
reg   [7:0]                            r_port_rxmac_down_regs            ;// �˿ڽ��շ���MAC�ر�ʹ��
reg   [7:0]                            r_port_broadcast_drop_regs        ;// �˿ڹ㲥֡����ʹ��
reg   [7:0]                            r_port_multicast_drop_regs        ;// �˿��鲥֡����ʹ��
reg   [7:0]                            r_port_loopback_drop_regs         ;// �˿ڻ���֡����ʹ��
reg   [7:0]                            r_port_force_recal_crc_regs       ;// �˿�ǿ�����¼���CRCʹ�� 
reg   [7:0]                            r_port_floodfrm_drop_regs         ;// �˿ڷ���֡����ʹ��   
reg   [7:0]                            r_port_multiflood_drop_regs       ;// �˿ڶಥ֡����ʹ�� 
reg   [7:0]                            r_port_acl_enable_regs                 ;// �˿� ACL ʹ��  


reg   [2:0]                            r_cfg_rxmac_port_sel              ;// �˿�ѡ��
reg   [47:0]                           r_port_mac_regs                   ;// �˿�1�� MAC ��ַ
reg                                    r_port_mac_vld_regs               ;// ʹ�ܶ˿� MAC ��ַ��Ч
reg   [10:0]                           r_port_mtu_regs                   ;// MTU����ֵ
reg   [PORT_NUM-1:0]                   r_port_mirror_frwd_regs           ;// ����ת���Ĵ���������Ӧ�Ķ˿���1���򱾶˿ڽ��յ����κ�ת������֡������ת��ֵ����1�Ķ˿�
reg   [15:0]                           r_port_flowctrl_cfg_regs          ;// ������������
reg   [4:0]                            r_port_rx_ultrashortinterval_num_0;// ֡���
reg   [4:0]                            r_port_rx_ultrashortinterval_num_1;// ֡���
reg   [4:0]                            r_port_rx_ultrashortinterval_num_2;// ֡���
reg   [4:0]                            r_port_rx_ultrashortinterval_num_3;// ֡���
reg   [4:0]                            r_port_rx_ultrashortinterval_num_4;// ֡���
reg   [4:0]                            r_port_rx_ultrashortinterval_num_5;// ֡���
reg   [4:0]                            r_port_rx_ultrashortinterval_num_6;// ֡���
reg   [4:0]                            r_port_rx_ultrashortinterval_num_7;// ֡���
/*========================================  ACL�Ĵ����źŶ��� ========================================*/

reg   [2:0]                            r_acl_port_sel                      ; // ѡ��Ҫ���õĶ˿�
reg                                    r_acl_clr_list_regs                 ; // ��ռĴ����б�
reg   [4:0]                            r_acl_item_sel_regs                 ; // ������Ŀѡ��
reg   [5:0]                            r_acl_item_waddr_regs               ; // ÿ����Ŀ���֧�ֱȶ� 64 �ֽ�
reg   [7:0]                            r_acl_item_din_regs                 ; // ��Ҫ�Ƚϵ��ֽ�����
reg                                    r_acl_item_we_regs                  ; // ����ʹ���ź�
reg   [15:0]                           r_acl_item_rslt_regs                ; // ƥ��Ľ��ֵ - [7:0] ���֡����, [15:8] ACLת��ָ���˿�
reg                                    r_acl_item_complete_regs            ; // �˿� ACL �����������ʹ���ź�
wire  [7:0]                            w_acl_list_rdy_regs                 ;

reg   [95:0]                           r_acl_item_dmac_code                ;
reg   [95:0]                           r_acl_item_smac_code                ;
reg   [63:0]                           r_acl_item_vlan_code                ;
reg   [31:0]                           r_acl_item_ethtype_code             ;
reg   [5:0]                            r_acl_item_action_pass_state        ;
reg   [15:0]                           r_acl_item_action_cb_streamhandle   ;
reg   [5:0]                            r_acl_item_action_flowctrl          ;
reg   [15:0]                           r_acl_item_action_txport            ;
/*--------------------------------------- Qbu_rx�Ĵ����źŶ��� ----------------------------------------*/
// �˿�0
reg                                    r_reset_0                           ;
reg                                    r_reset_1                           ;
reg                                    r_reset_2                           ;
reg                                    r_reset_3                           ;
reg                                    r_reset_4                           ;
reg                                    r_reset_5                           ;
reg                                    r_reset_6                           ;
reg                                    r_reset_7                           ;

/*========================================  ͨ�üĴ��������źŹ��� ========================================*/
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_refresh_list_pulse        <= 1'b0;
        r_switch_err_cnt_clr        <= 1'b0;
        r_switch_err_cnt_stat       <= 1'b0;
    end else begin
        r_refresh_list_pulse        <= i_refresh_list_pulse;
        r_switch_err_cnt_clr        <= i_switch_err_cnt_clr;
        r_switch_err_cnt_stat       <= i_switch_err_cnt_stat;
    end
end
/*========================================  �Ĵ�����д�����źŹ��� ========================================*/
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_reg_bus_we          <= 1'b0;
        r_reg_bus_addr        <= {REG_ADDR_BUS_WIDTH{1'b0}};
        r_reg_bus_data        <= {REG_DATA_BUS_WIDTH{1'b0}};
        r_reg_bus_data_vld    <= 1'b0;
        r_reg_bus_re          <= 1'b0;
        r_reg_bus_raddr       <= {REG_ADDR_BUS_WIDTH{1'b0}};
    end else begin
        r_reg_bus_we          <= i_switch_reg_bus_we;
        r_reg_bus_addr        <= i_switch_reg_bus_we_addr;
        r_reg_bus_data        <= i_switch_reg_bus_we_din;
        r_reg_bus_data_vld    <= i_switch_reg_bus_we_din_v;
        r_reg_bus_re          <= i_switch_reg_bus_rd;
        r_reg_bus_raddr       <= i_switch_reg_bus_rd_addr;
    end
end

always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
		r_hash_ploy_regs <= 16'h180F;
        r_hash_init_val_regs <= 16'hFFFF;
        r_hash_regs_vld <= 1'b0;
        r_port_rxmac_down_regs <= 8'hFF;
        r_port_acl_enable_regs <= 8'hFF;
        r_port_broadcast_drop_regs <= 8'b0;
        r_port_multicast_drop_regs <= 8'b0;
        r_port_loopback_drop_regs <= 8'hFF;
        r_port_force_recal_crc_regs <= 8'b0;
        r_port_floodfrm_drop_regs <= 8'b1;
        r_port_multiflood_drop_regs <= 8'b0;
        r_cfg_rxmac_port_sel <= 3'b0;
        r_port_mac_regs <= 48'b0;
        r_port_mac_vld_regs <= 1'b0;
        r_port_mtu_regs <= 11'd1600;
        r_port_mirror_frwd_regs <= 8'b0;
        r_port_flowctrl_cfg_regs <= 16'b0;
        //r_port_rx_ultrashortinterval_num <= 5'd31;
    end else begin
        r_hash_ploy_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_HASH_PLOY ? r_reg_bus_data[15:0] : r_hash_ploy_regs;
        r_hash_init_val_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_HASH_INIT_VAL ? r_reg_bus_data[15:0] : r_hash_init_val_regs;
        r_hash_regs_vld <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_HASH_INIT_VAL ? 1'b1 : 1'b0;
        r_port_rxmac_down_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_RXMAC_DOWN ? r_reg_bus_data[7:0] : r_port_rxmac_down_regs;
        r_port_broadcast_drop_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_BROADCAST_DROP ? r_reg_bus_data[7:0] : r_port_broadcast_drop_regs;
        r_port_multicast_drop_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_MULTICAST_DROP ? r_reg_bus_data[7:0] : r_port_multicast_drop_regs;
        r_port_loopback_drop_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_LOOKBACK_DROP ? r_reg_bus_data[7:0] : r_port_loopback_drop_regs;
        r_port_force_recal_crc_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_FORCE_RECAL_CRC ? r_reg_bus_data[7:0] : r_port_force_recal_crc_regs;
        r_port_floodfrm_drop_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_FLOODFRM_DROP ? r_reg_bus_data[7:0] : r_port_floodfrm_drop_regs;
        r_port_multiflood_drop_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_MULTIFLOOD_DROP ? r_reg_bus_data[7:0] : r_port_multiflood_drop_regs;
        r_cfg_rxmac_port_sel <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_CFG_RXMAC_PORT_SEL ? r_reg_bus_data[2:0] : r_cfg_rxmac_port_sel;
        r_port_mac_regs[47:32] <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORTMAC0 ? r_reg_bus_data[15:0] : r_port_mac_regs[47:32];
        r_port_mac_regs[31:16] <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORTMAC1 ? r_reg_bus_data[15:0] : r_port_mac_regs[31:16];
        r_port_mac_regs[15:0] <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORTMAC2 ? r_reg_bus_data[15:0] : r_port_mac_regs[15:0];
        r_port_mac_vld_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORTMAC_VALID ? r_reg_bus_data[0] : r_port_mac_vld_regs;
        r_port_mtu_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORTMTU ? r_reg_bus_data[10:0] : r_port_mtu_regs;
        r_port_mirror_frwd_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_MIRROR_FRWD ? r_reg_bus_data[7:0] : r_port_mirror_frwd_regs;
        r_port_flowctrl_cfg_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_FLOWCTRL_CFG ? r_reg_bus_data[15:0] : r_port_flowctrl_cfg_regs;
        //r_port_rx_ultrashortinterval_num <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_RX_ULTRASHORTINTERVAL_NUM ? r_reg_bus_data[4:0] : r_port_rx_ultrashortinterval_num;
        r_port_acl_enable_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_ACL_ENABLE ? r_reg_bus_data[7:0] : r_port_acl_enable_regs;
    end
end
// �˿�1
assign o_hash_ploy_regs_0 = r_hash_ploy_regs;
assign o_hash_init_val_regs_0 = r_hash_init_val_regs;
assign o_hash_regs_vld_0 = r_hash_regs_vld;
assign o_port_rxmac_down_regs_0 = r_port_rxmac_down_regs[0];
assign o_port_broadcast_drop_regs_0 = r_port_broadcast_drop_regs[0];
assign o_port_multicast_drop_regs_0 = r_port_multicast_drop_regs[0];
assign o_port_loopback_drop_regs_0 = r_port_loopback_drop_regs[0];
assign o_port_mac_regs_0 = r_cfg_rxmac_port_sel == 3'b000 ? r_port_mac_regs[47:0] : 48'b0;
assign o_port_mac_vld_regs_0 = r_cfg_rxmac_port_sel == 3'b000 ? r_port_mac_vld_regs : 1'b0;
assign o_port_mtu_regs_0 = r_cfg_rxmac_port_sel == 3'b000 ? r_port_mtu_regs : 8'b0;
assign o_port_mirror_frwd_regs_0 = r_cfg_rxmac_port_sel == 3'b000 ? r_port_mirror_frwd_regs : 8'b0;
assign o_port_flowctrl_cfg_regs_0 = r_cfg_rxmac_port_sel == 3'b000 ? r_port_flowctrl_cfg_regs : 16'b0;
//assign o_port_rx_ultrashortinterval_num_0 = r_cfg_rxmac_port_sel == 3'b000 ? r_port_rx_ultrashortinterval_num : 5'b0;

// �˿�2
assign o_hash_ploy_regs_1 = r_hash_ploy_regs;
assign o_hash_init_val_regs_1 = r_hash_init_val_regs;
assign o_hash_regs_vld_1 = r_hash_regs_vld;
assign o_port_rxmac_down_regs_1 = r_port_rxmac_down_regs[1];
assign o_port_broadcast_drop_regs_1 = r_port_broadcast_drop_regs[1];
assign o_port_multicast_drop_regs_1 = r_port_multicast_drop_regs[1];
assign o_port_loopback_drop_regs_1 = r_port_loopback_drop_regs[1];
assign o_port_mac_regs_1 = r_cfg_rxmac_port_sel == 3'b001 ? r_port_mac_regs[47:0] : 48'b0;
assign o_port_mac_vld_regs_1 = r_cfg_rxmac_port_sel == 3'b001 ? r_port_mac_vld_regs : 1'b0;
assign o_port_mtu_regs_1 = r_cfg_rxmac_port_sel == 3'b001 ? r_port_mtu_regs : 8'b0;
assign o_port_mirror_frwd_regs_1 = r_cfg_rxmac_port_sel == 3'b001 ? r_port_mirror_frwd_regs : 8'b0;
assign o_port_flowctrl_cfg_regs_1 = r_cfg_rxmac_port_sel == 3'b001 ? r_port_flowctrl_cfg_regs : 16'b0;
//assign o_port_rx_ultrashortinterval_num_1 = r_cfg_rxmac_port_sel == 3'b001 ? r_port_rx_ultrashortinterval_num : 5'b0;

// �˿�3
assign o_hash_ploy_regs_2 = r_hash_ploy_regs;
assign o_hash_init_val_regs_2 = r_hash_init_val_regs;
assign o_hash_regs_vld_2 = r_hash_regs_vld;
assign o_port_rxmac_down_regs_2 = r_port_rxmac_down_regs[2];
assign o_port_broadcast_drop_regs_2 = r_port_broadcast_drop_regs[2];
assign o_port_multicast_drop_regs_2 = r_port_multicast_drop_regs[2];
assign o_port_loopback_drop_regs_2 = r_port_loopback_drop_regs[2];
assign o_port_mac_regs_2 = r_cfg_rxmac_port_sel == 3'b010 ? r_port_mac_regs[47:0] : 48'b0;
assign o_port_mac_vld_regs_2 = r_cfg_rxmac_port_sel == 3'b010 ? r_port_mac_vld_regs : 1'b0;
assign o_port_mtu_regs_2 = r_cfg_rxmac_port_sel == 3'b010 ? r_port_mtu_regs : 8'b0;
assign o_port_mirror_frwd_regs_2 = r_cfg_rxmac_port_sel == 3'b010 ? r_port_mirror_frwd_regs : 8'b0;
assign o_port_flowctrl_cfg_regs_2 = r_cfg_rxmac_port_sel == 3'b010 ? r_port_flowctrl_cfg_regs : 16'b0;
//assign o_port_rx_ultrashortinterval_num_2 = r_cfg_rxmac_port_sel == 3'b010 ? r_port_rx_ultrashortinterval_num : 5'b0;

// �˿�4
assign o_hash_ploy_regs_3 = r_hash_ploy_regs;
assign o_hash_init_val_regs_3 = r_hash_init_val_regs;
assign o_hash_regs_vld_3 = r_hash_regs_vld;
assign o_port_rxmac_down_regs_3 = r_port_rxmac_down_regs[3];
assign o_port_broadcast_drop_regs_3 = r_port_broadcast_drop_regs[3];
assign o_port_multicast_drop_regs_3 = r_port_multicast_drop_regs[3];
assign o_port_loopback_drop_regs_3 = r_port_loopback_drop_regs[3];
assign o_port_mac_regs_3 = r_cfg_rxmac_port_sel == 3'b011 ? r_port_mac_regs[47:0] : 48'b0;
assign o_port_mac_vld_regs_3 = r_cfg_rxmac_port_sel == 3'b011 ? r_port_mac_vld_regs : 1'b0;
assign o_port_mtu_regs_3 = r_cfg_rxmac_port_sel == 3'b011 ? r_port_mtu_regs : 8'b0;
assign o_port_mirror_frwd_regs_3 = r_cfg_rxmac_port_sel == 3'b011 ? r_port_mirror_frwd_regs : 8'b0;
assign o_port_flowctrl_cfg_regs_3 = r_cfg_rxmac_port_sel == 3'b011 ? r_port_flowctrl_cfg_regs : 16'b0;
//assign o_port_rx_ultrashortinterval_num_3 = r_cfg_rxmac_port_sel == 3'b011 ? r_port_rx_ultrashortinterval_num : 5'b0;

// �˿�5
assign o_hash_ploy_regs_4 = r_hash_ploy_regs;
assign o_hash_init_val_regs_4 = r_hash_init_val_regs;
assign o_hash_regs_vld_4 = r_hash_regs_vld;
assign o_port_rxmac_down_regs_4 = r_port_rxmac_down_regs[4];
assign o_port_broadcast_drop_regs_4 = r_port_broadcast_drop_regs[4];
assign o_port_multicast_drop_regs_4 = r_port_multicast_drop_regs[4];
assign o_port_loopback_drop_regs_4 = r_port_loopback_drop_regs[4];
assign o_port_mac_regs_4 = r_cfg_rxmac_port_sel == 3'b100 ? r_port_mac_regs[47:0] : 48'b0;
assign o_port_mac_vld_regs_4 = r_cfg_rxmac_port_sel == 3'b100 ? r_port_mac_vld_regs : 1'b0;
assign o_port_mtu_regs_4 = r_cfg_rxmac_port_sel == 3'b100 ? r_port_mtu_regs : 8'b0;
assign o_port_mirror_frwd_regs_4 = r_cfg_rxmac_port_sel == 3'b100 ? r_port_mirror_frwd_regs : 8'b0;
assign o_port_flowctrl_cfg_regs_4 = r_cfg_rxmac_port_sel == 3'b100 ? r_port_flowctrl_cfg_regs : 16'b0;
//assign o_port_rx_ultrashortinterval_num_4 = r_cfg_rxmac_port_sel == 3'b100 ? r_port_rx_ultrashortinterval_num : 5'b0;

// �˿�6
assign o_hash_ploy_regs_5 = r_hash_ploy_regs;
assign o_hash_init_val_regs_5 = r_hash_init_val_regs;
assign o_hash_regs_vld_5 = r_hash_regs_vld;
assign o_port_rxmac_down_regs_5 = r_port_rxmac_down_regs[5];
assign o_port_broadcast_drop_regs_5 = r_port_broadcast_drop_regs[5];
assign o_port_multicast_drop_regs_5 = r_port_multicast_drop_regs[5];
assign o_port_loopback_drop_regs_5 = r_port_loopback_drop_regs[5];
assign o_port_mac_regs_5 = r_cfg_rxmac_port_sel == 3'b101 ? r_port_mac_regs[47:0] : 48'b0;
assign o_port_mac_vld_regs_5 = r_cfg_rxmac_port_sel == 3'b101 ? r_port_mac_vld_regs : 1'b0;
assign o_port_mtu_regs_5 = r_cfg_rxmac_port_sel == 3'b101 ? r_port_mtu_regs : 8'b0;
assign o_port_mirror_frwd_regs_5 = r_cfg_rxmac_port_sel == 3'b101 ? r_port_mirror_frwd_regs : 8'b0;
assign o_port_flowctrl_cfg_regs_5 = r_cfg_rxmac_port_sel == 3'b101 ? r_port_flowctrl_cfg_regs : 16'b0;
//assign o_port_rx_ultrashortinterval_num_5 = r_cfg_rxmac_port_sel == 3'b101 ? r_port_rx_ultrashortinterval_num : 5'b0;

// �˿�7
assign o_hash_ploy_regs_6 = r_hash_ploy_regs;
assign o_hash_init_val_regs_6 = r_hash_init_val_regs;
assign o_hash_regs_vld_6 = r_hash_regs_vld;
assign o_port_rxmac_down_regs_6 = r_port_rxmac_down_regs[6];
assign o_port_broadcast_drop_regs_6 = r_port_broadcast_drop_regs[6];
assign o_port_multicast_drop_regs_6 = r_port_multicast_drop_regs[6];
assign o_port_loopback_drop_regs_6 = r_port_loopback_drop_regs[6];
assign o_port_mac_regs_6 = r_cfg_rxmac_port_sel == 3'b110 ? r_port_mac_regs[47:0] : 48'b0;
assign o_port_mac_vld_regs_6 = r_cfg_rxmac_port_sel == 3'b110 ? r_port_mac_vld_regs : 1'b0;
assign o_port_mtu_regs_6 = r_cfg_rxmac_port_sel == 3'b110 ? r_port_mtu_regs : 8'b0;
assign o_port_mirror_frwd_regs_6 = r_cfg_rxmac_port_sel == 3'b110 ? r_port_mirror_frwd_regs : 8'b0;
assign o_port_flowctrl_cfg_regs_6 = r_cfg_rxmac_port_sel == 3'b110 ? r_port_flowctrl_cfg_regs : 16'b0;
//assign o_port_rx_ultrashortinterval_num_6 = r_cfg_rxmac_port_sel == 3'b110 ? r_port_rx_ultrashortinterval_num : 5'b0;

// �˿�8
assign o_hash_ploy_regs_7 = r_hash_ploy_regs;
assign o_hash_init_val_regs_7 = r_hash_init_val_regs;
assign o_hash_regs_vld_7 = r_hash_regs_vld;
assign o_port_rxmac_down_regs_7 = r_port_rxmac_down_regs[7];
assign o_port_broadcast_drop_regs_7 = r_port_broadcast_drop_regs[7];
assign o_port_multicast_drop_regs_7 = r_port_multicast_drop_regs[7];
assign o_port_loopback_drop_regs_7 = r_port_loopback_drop_regs[7];
assign o_port_mac_regs_7 = r_cfg_rxmac_port_sel == 3'b111 ? r_port_mac_regs[47:0] : 48'b0;
assign o_port_mac_vld_regs_7 = r_cfg_rxmac_port_sel == 3'b111 ? r_port_mac_vld_regs : 1'b0;
assign o_port_mtu_regs_7 = r_cfg_rxmac_port_sel == 3'b111 ? r_port_mtu_regs : 8'b0;
assign o_port_mirror_frwd_regs_7 = r_cfg_rxmac_port_sel == 3'b111 ? r_port_mirror_frwd_regs : 8'b0;
assign o_port_flowctrl_cfg_regs_7 = r_cfg_rxmac_port_sel == 3'b111 ? r_port_flowctrl_cfg_regs : 16'b0;
//assign o_port_rx_ultrashortinterval_num_7 = r_cfg_rxmac_port_sel == 3'b111 ? r_port_rx_ultrashortinterval_num : 5'b0;

always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_port_rx_ultrashortinterval_num_0 <= 5'd31;
        r_port_rx_ultrashortinterval_num_1 <= 5'd31;
        r_port_rx_ultrashortinterval_num_2 <= 5'd31;
        r_port_rx_ultrashortinterval_num_3 <= 5'd31;
        r_port_rx_ultrashortinterval_num_4 <= 5'd31;
        r_port_rx_ultrashortinterval_num_5 <= 5'd31;
        r_port_rx_ultrashortinterval_num_6 <= 5'd31;
        r_port_rx_ultrashortinterval_num_7 <= 5'd31;
    end else begin
        r_port_rx_ultrashortinterval_num_0 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_RX_ULTRASHORTINTERVAL_NUM_0 ? r_reg_bus_data[4:0] : r_port_rx_ultrashortinterval_num_0;
        r_port_rx_ultrashortinterval_num_1 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_RX_ULTRASHORTINTERVAL_NUM_1 ? r_reg_bus_data[4:0] : r_port_rx_ultrashortinterval_num_1;
        r_port_rx_ultrashortinterval_num_2 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_RX_ULTRASHORTINTERVAL_NUM_2 ? r_reg_bus_data[4:0] : r_port_rx_ultrashortinterval_num_2;
        r_port_rx_ultrashortinterval_num_3 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_RX_ULTRASHORTINTERVAL_NUM_3 ? r_reg_bus_data[4:0] : r_port_rx_ultrashortinterval_num_3;
        r_port_rx_ultrashortinterval_num_4 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_RX_ULTRASHORTINTERVAL_NUM_4 ? r_reg_bus_data[4:0] : r_port_rx_ultrashortinterval_num_4;
        r_port_rx_ultrashortinterval_num_5 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_RX_ULTRASHORTINTERVAL_NUM_5 ? r_reg_bus_data[4:0] : r_port_rx_ultrashortinterval_num_5;
        r_port_rx_ultrashortinterval_num_6 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_RX_ULTRASHORTINTERVAL_NUM_6 ? r_reg_bus_data[4:0] : r_port_rx_ultrashortinterval_num_6;
        r_port_rx_ultrashortinterval_num_7 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_PORT_RX_ULTRASHORTINTERVAL_NUM_7 ? r_reg_bus_data[4:0] : r_port_rx_ultrashortinterval_num_7;
    end
end

assign o_port_rx_ultrashortinterval_num_0 = r_port_rx_ultrashortinterval_num_0;
assign o_port_rx_ultrashortinterval_num_1 = r_port_rx_ultrashortinterval_num_1;
assign o_port_rx_ultrashortinterval_num_2 = r_port_rx_ultrashortinterval_num_2;
assign o_port_rx_ultrashortinterval_num_3 = r_port_rx_ultrashortinterval_num_3;
assign o_port_rx_ultrashortinterval_num_4 = r_port_rx_ultrashortinterval_num_4;
assign o_port_rx_ultrashortinterval_num_5 = r_port_rx_ultrashortinterval_num_5;
assign o_port_rx_ultrashortinterval_num_6 = r_port_rx_ultrashortinterval_num_6;
assign o_port_rx_ultrashortinterval_num_7 = r_port_rx_ultrashortinterval_num_7;

/*========================================  ACL�Ĵ���д�����źŹ��� ========================================*/

always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_acl_port_sel <= 3'b0;
        r_acl_clr_list_regs <= 1'b0;
        r_acl_item_sel_regs <= 5'b0;
    end else begin
        r_acl_port_sel <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_CFG_ACL_PORT_SEL ? r_reg_bus_data[2:0] : r_acl_port_sel;
        r_acl_clr_list_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_CFG_ACL_CLR_LIST ? r_reg_bus_data[0] : r_acl_clr_list_regs;
        r_acl_item_sel_regs <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_CFG_ACL_ITEM_SEL ? r_reg_bus_data[4:0] : r_acl_item_sel_regs;
    end
end

// ACL��Ŀ����д����
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_acl_item_dmac_code <= 96'b0;
        r_acl_item_smac_code <= 96'b0;
        r_acl_item_vlan_code <= 64'b0;
        r_acl_item_ethtype_code <= 32'b0;
        r_acl_item_action_pass_state <= 6'b0;
        r_acl_item_action_cb_streamhandle <= 16'b0;
        r_acl_item_action_flowctrl <= 6'b0;
        r_acl_item_action_txport <= 16'b0;
    end else begin
        if (r_reg_bus_we && r_reg_bus_data_vld) begin
            case (r_reg_bus_addr)
                REG_CFG_ACL_ITEM_DMAC_CODE_1: r_acl_item_dmac_code[15:0]  <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_DMAC_CODE_2: r_acl_item_dmac_code[31:16] <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_DMAC_CODE_3: r_acl_item_dmac_code[47:32] <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_DMAC_CODE_4: r_acl_item_dmac_code[63:48] <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_DMAC_CODE_5: r_acl_item_dmac_code[79:64] <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_DMAC_CODE_6: r_acl_item_dmac_code[95:80] <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_SMAC_CODE_1: r_acl_item_smac_code[15:0]  <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_SMAC_CODE_2: r_acl_item_smac_code[31:16] <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_SMAC_CODE_3: r_acl_item_smac_code[47:32] <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_SMAC_CODE_4: r_acl_item_smac_code[63:48] <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_SMAC_CODE_5: r_acl_item_smac_code[79:64] <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_SMAC_CODE_6: r_acl_item_smac_code[95:80] <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_VLAN_CODE_1: r_acl_item_vlan_code[15:0]  <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_VLAN_CODE_2: r_acl_item_vlan_code[31:16] <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_VLAN_CODE_3: r_acl_item_vlan_code[47:32] <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_VLAN_CODE_4: r_acl_item_vlan_code[63:48] <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_ETHTYPE_CODE_1: r_acl_item_ethtype_code[15:0] <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_ETHTYPE_CODE_2: r_acl_item_ethtype_code[31:16] <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_ACTION_PASS_STATE: r_acl_item_action_pass_state <= r_reg_bus_data[5:0];
                REG_CFG_ACL_ITEM_ACTION_CB_STREAMHANDLE: r_acl_item_action_cb_streamhandle <= r_reg_bus_data[15:0];
                REG_CFG_ACL_ITEM_ACTION_FLOWCTRL: r_acl_item_action_flowctrl <= r_reg_bus_data[5:0];
                REG_CFG_ACL_ITEM_ACTION_TXPORT: r_acl_item_action_txport <= r_reg_bus_data[15:0];
            endcase
        end
    end
end


// �˿�1
assign o_acl_clr_list_regs_0 = r_acl_port_sel == 3'b000 ? r_acl_clr_list_regs : 1'b0;
assign o_acl_item_sel_regs_0 = r_acl_port_sel == 3'b000 ? r_acl_item_sel_regs : 5'b0;
// �˿�2
assign o_acl_clr_list_regs_1 = r_acl_port_sel == 3'b001 ? r_acl_clr_list_regs : 1'b0;
assign o_acl_item_sel_regs_1 = r_acl_port_sel == 3'b001 ? r_acl_item_sel_regs : 5'b0;
// �˿�3
assign o_acl_clr_list_regs_2 = r_acl_port_sel == 3'b010 ? r_acl_clr_list_regs : 1'b0;
assign o_acl_item_sel_regs_2 = r_acl_port_sel == 3'b010 ? r_acl_item_sel_regs : 5'b0;
// �˿�4
assign o_acl_clr_list_regs_3 = r_acl_port_sel == 3'b011 ? r_acl_clr_list_regs : 1'b0;
assign o_acl_item_sel_regs_3 = r_acl_port_sel == 3'b011 ? r_acl_item_sel_regs : 5'b0;
// �˿�5
assign o_acl_clr_list_regs_4 = r_acl_port_sel == 3'b100 ? r_acl_clr_list_regs : 1'b0;
assign o_acl_item_sel_regs_4 = r_acl_port_sel == 3'b100 ? r_acl_item_sel_regs : 5'b0;
// �˿�6
assign o_acl_clr_list_regs_5 = r_acl_port_sel == 3'b101 ? r_acl_clr_list_regs : 1'b0;
assign o_acl_item_sel_regs_5 = r_acl_port_sel == 3'b101 ? r_acl_item_sel_regs : 5'b0;
// �˿�7
assign o_acl_clr_list_regs_6 = r_acl_port_sel == 3'b110 ? r_acl_clr_list_regs : 1'b0;
assign o_acl_item_sel_regs_6 = r_acl_port_sel == 3'b110 ? r_acl_item_sel_regs : 5'b0;
// �˿�8
assign o_acl_clr_list_regs_7 = r_acl_port_sel == 3'b111 ? r_acl_clr_list_regs : 1'b0;
assign o_acl_item_sel_regs_7 = r_acl_port_sel == 3'b111 ? r_acl_item_sel_regs : 5'b0;

/*========================================  qbu_rx�Ĵ���д�����źŹ��� ========================================*/

// QBU��λ�Ĵ���д���� - ���ж˿�
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_reset_0 <= 1'b0;
        r_reset_1 <= 1'b0;
        r_reset_2 <= 1'b0;
        r_reset_3 <= 1'b0;
        r_reset_4 <= 1'b0;
        r_reset_5 <= 1'b0;
        r_reset_6 <= 1'b0;
        r_reset_7 <= 1'b0;
    end else begin
        r_reset_0 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_QBU_RESET_0 ? r_reg_bus_data[0] : 1'b0;
        r_reset_1 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_QBU_RESET_1 ? r_reg_bus_data[0] : 1'b0;
        r_reset_2 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_QBU_RESET_2 ? r_reg_bus_data[0] : 1'b0;
        r_reset_3 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_QBU_RESET_3 ? r_reg_bus_data[0] : 1'b0;
        r_reset_4 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_QBU_RESET_4 ? r_reg_bus_data[0] : 1'b0;
        r_reset_5 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_QBU_RESET_5 ? r_reg_bus_data[0] : 1'b0;
        r_reset_6 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_QBU_RESET_6 ? r_reg_bus_data[0] : 1'b0;
        r_reset_7 <= r_reg_bus_we == 1'b1 && r_reg_bus_data_vld == 1'b1 && r_reg_bus_addr == REG_QBU_RESET_7 ? r_reg_bus_data[0] : 1'b0;
    end
end

assign o_reset_0 = r_reset_0;
assign o_reset_1 = r_reset_1;
assign o_reset_2 = r_reset_2;
assign o_reset_3 = r_reset_3;
assign o_reset_4 = r_reset_4;
assign o_reset_5 = r_reset_5;
assign o_reset_6 = r_reset_6;
assign o_reset_7 = r_reset_7;

assign w_acl_list_rdy_regs = {i_acl_list_rdy_regs_7,i_acl_list_rdy_regs_6,i_acl_list_rdy_regs_5,i_acl_list_rdy_regs_4,
                              i_acl_list_rdy_regs_3,i_acl_list_rdy_regs_2,i_acl_list_rdy_regs_1,i_acl_list_rdy_regs_0};
/*========================================= �Ĵ����������߼� =========================================*/
// �Ĵ����������߼�
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_reg_bus_rdata <= {REG_DATA_BUS_WIDTH{1'b0}};
    end else if (r_reg_bus_re) begin
        case (r_reg_bus_raddr)
            // rxmac ͨ��
            REG_HASH_PLOY:    r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_hash_ploy_regs; 
            REG_HASH_INIT_VAL:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_hash_init_val_regs; 
            REG_PORT_RXMAC_DOWN:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_port_rxmac_down_regs; 
            REG_PORT_ACL_ENABLE:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_port_acl_enable_regs; 
            REG_PORT_BROADCAST_DROP:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_port_broadcast_drop_regs; 
            REG_PORT_MULTICAST_DROP:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_port_multicast_drop_regs; 
            REG_PORT_LOOKBACK_DROP:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_port_loopback_drop_regs; 
            REG_PORT_FORCE_RECAL_CRC:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_port_force_recal_crc_regs; 
            REG_PORT_FLOODFRM_DROP:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_port_floodfrm_drop_regs; 
            REG_PORT_MULTIFLOOD_DROP:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_port_multiflood_drop_regs; 
            REG_CFG_RXMAC_PORT_SEL:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_cfg_rxmac_port_sel; 
            REG_PORTMTU:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_port_mtu_regs; 
            REG_PORTMAC0:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_port_mac_regs[47:32]; 
            REG_PORTMAC1:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_port_mac_regs[31:16];
            REG_PORTMAC2:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_port_mac_regs[15:0];
            REG_PORTMAC_VALID:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_port_mac_vld_regs;
            REG_PORT_MIRROR_FRWD:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_port_mirror_frwd_regs;
            REG_PORT_FLOWCTRL_CFG:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_port_flowctrl_cfg_regs;
            // acl�Ĵ���
            REG_CFG_ACL_PORT_SEL:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_port_sel;
            REG_CFG_ACL_CLR_LIST:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_clr_list_regs;
            REG_CFG_ACL_LIST_RDY:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | w_acl_list_rdy_regs;
            REG_CFG_ACL_ITEM_SEL:  r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_sel_regs;
            REG_CFG_ACL_ITEM_DMAC_CODE_1: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_dmac_code[15:0];
            REG_CFG_ACL_ITEM_DMAC_CODE_2: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_dmac_code[31:16];
            REG_CFG_ACL_ITEM_DMAC_CODE_3: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_dmac_code[47:32];
            REG_CFG_ACL_ITEM_DMAC_CODE_4: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_dmac_code[63:48];
            REG_CFG_ACL_ITEM_DMAC_CODE_5: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_dmac_code[79:64];
            REG_CFG_ACL_ITEM_DMAC_CODE_6: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_dmac_code[95:80];
            REG_CFG_ACL_ITEM_SMAC_CODE_1: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_smac_code[15:0];
            REG_CFG_ACL_ITEM_SMAC_CODE_2: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_smac_code[31:16];
            REG_CFG_ACL_ITEM_SMAC_CODE_3: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_smac_code[47:32];
            REG_CFG_ACL_ITEM_SMAC_CODE_4: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_smac_code[63:48];
            REG_CFG_ACL_ITEM_SMAC_CODE_5: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_smac_code[79:64];
            REG_CFG_ACL_ITEM_SMAC_CODE_6: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_smac_code[95:80];
            REG_CFG_ACL_ITEM_VLAN_CODE_1: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_vlan_code[15:0];
            REG_CFG_ACL_ITEM_VLAN_CODE_2: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_vlan_code[31:16];
            REG_CFG_ACL_ITEM_VLAN_CODE_3: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_vlan_code[47:32];
            REG_CFG_ACL_ITEM_VLAN_CODE_4: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_vlan_code[63:48];
            REG_CFG_ACL_ITEM_ETHTYPE_CODE_1: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_ethtype_code[15:0];
            REG_CFG_ACL_ITEM_ETHTYPE_CODE_2: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_ethtype_code[31:16];
            REG_CFG_ACL_ITEM_ACTION_PASS_STATE: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_action_pass_state;
            REG_CFG_ACL_ITEM_ACTION_CB_STREAMHANDLE: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_action_cb_streamhandle;
            REG_CFG_ACL_ITEM_ACTION_FLOWCTRL: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_action_flowctrl;
            REG_CFG_ACL_ITEM_ACTION_TXPORT: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | r_acl_item_action_txport;
            // rxmac port
            // �˿�1
            REG_PORT_RX_BYTE_CNT_0:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_byte_cnt_0;
            REG_PORT_RX_FRAME_CNT_0:    r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_frame_cnt_0;
            REG_PORT_DIAG_STATE_0:      r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, i_port_diag_state_0};
            //REG_PORT_RX_ULTRASHORT_FRM_CNT_0: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_ultrashort_frm_cnt_0; 
            //REG_PORT_RX_OVERLENGTH_FRM_CNT_0: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_overlength_frm_cnt_0; 
            //REG_PORT_RX_CRCERR_FRM_CNT_0: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_crcerr_frm_cnt_0;     
            //REG_PORT_RX_LOOKBACK_FRM_CNT_0: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_lookback_frm_cnt_0; 
            REG_PORT_BROADFLOW_DROP_CNT_0: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_broadflow_drop_cnt_0; 
            REG_PORT_MULTIFLOW_DROP_CNT_0: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_multiflow_drop_cnt_0; 
            // �˿�2
            REG_PORT_RX_BYTE_CNT_1:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_byte_cnt_1;
            REG_PORT_RX_FRAME_CNT_1:    r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_frame_cnt_1;
            REG_PORT_DIAG_STATE_1:      r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, i_port_diag_state_1};
            //REG_PORT_RX_ULTRASHORT_FRM_CNT_1: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_ultrashort_frm_cnt_1; 
            //REG_PORT_RX_OVERLENGTH_FRM_CNT_1: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_overlength_frm_cnt_1; 
            //REG_PORT_RX_CRCERR_FRM_CNT_1: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_crcerr_frm_cnt_1;     
            //REG_PORT_RX_LOOKBACK_FRM_CNT_1: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_lookback_frm_cnt_1; 
            REG_PORT_BROADFLOW_DROP_CNT_1: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_broadflow_drop_cnt_1; 
            REG_PORT_MULTIFLOW_DROP_CNT_1: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_multiflow_drop_cnt_1; 
            // �˿�3
            REG_PORT_RX_BYTE_CNT_2:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_byte_cnt_2;
            REG_PORT_RX_FRAME_CNT_2:    r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_frame_cnt_2;
            REG_PORT_DIAG_STATE_2:      r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, i_port_diag_state_2};
            //REG_PORT_RX_ULTRASHORT_FRM_CNT_2: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_ultrashort_frm_cnt_2; 
            //REG_PORT_RX_OVERLENGTH_FRM_CNT_2: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_overlength_frm_cnt_2; 
            //REG_PORT_RX_CRCERR_FRM_CNT_2: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_crcerr_frm_cnt_2;     
            //REG_PORT_RX_LOOKBACK_FRM_CNT_2: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_lookback_frm_cnt_2; 
            REG_PORT_BROADFLOW_DROP_CNT_2: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_broadflow_drop_cnt_2; 
            REG_PORT_MULTIFLOW_DROP_CNT_2: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_multiflow_drop_cnt_2; 
            // �˿�4
            REG_PORT_RX_BYTE_CNT_3:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_byte_cnt_3;
            REG_PORT_RX_FRAME_CNT_3:    r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_frame_cnt_3;
            REG_PORT_DIAG_STATE_3:      r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, i_port_diag_state_3};
            //REG_PORT_RX_ULTRASHORT_FRM_CNT_3: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_ultrashort_frm_cnt_3; 
            //REG_PORT_RX_OVERLENGTH_FRM_CNT_3: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_overlength_frm_cnt_3; 
            //REG_PORT_RX_CRCERR_FRM_CNT_3: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_crcerr_frm_cnt_3;     
            //REG_PORT_RX_LOOKBACK_FRM_CNT_3: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_lookback_frm_cnt_3; 
            REG_PORT_BROADFLOW_DROP_CNT_3: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_broadflow_drop_cnt_3; 
            REG_PORT_MULTIFLOW_DROP_CNT_3: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_multiflow_drop_cnt_3; 
            // �˿�5
            REG_PORT_RX_BYTE_CNT_4:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_byte_cnt_4;
            REG_PORT_RX_FRAME_CNT_4:    r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_frame_cnt_4;
            REG_PORT_DIAG_STATE_4:      r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, i_port_diag_state_4};
            //REG_PORT_RX_ULTRASHORT_FRM_CNT_4: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_ultrashort_frm_cnt_4; 
            //REG_PORT_RX_OVERLENGTH_FRM_CNT_4: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_overlength_frm_cnt_4; 
            //REG_PORT_RX_CRCERR_FRM_CNT_4: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_crcerr_frm_cnt_4;     
            //REG_PORT_RX_LOOKBACK_FRM_CNT_4: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_lookback_frm_cnt_4; 
            REG_PORT_BROADFLOW_DROP_CNT_4: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_broadflow_drop_cnt_4; 
            REG_PORT_MULTIFLOW_DROP_CNT_4: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_multiflow_drop_cnt_4; 
            // �˿�6
            REG_PORT_RX_BYTE_CNT_5:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_byte_cnt_5;
            REG_PORT_RX_FRAME_CNT_5:    r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_frame_cnt_5;
            REG_PORT_DIAG_STATE_5:      r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, i_port_diag_state_5};
            //REG_PORT_RX_ULTRASHORT_FRM_CNT_5: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_ultrashort_frm_cnt_5; 
            //REG_PORT_RX_OVERLENGTH_FRM_CNT_5: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_overlength_frm_cnt_5; 
            //REG_PORT_RX_CRCERR_FRM_CNT_5: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_crcerr_frm_cnt_5;     
            //REG_PORT_RX_LOOKBACK_FRM_CNT_5: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_lookback_frm_cnt_5; 
            REG_PORT_BROADFLOW_DROP_CNT_5: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_broadflow_drop_cnt_5; 
            REG_PORT_MULTIFLOW_DROP_CNT_5: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_multiflow_drop_cnt_5; 
            // �˿�7
            REG_PORT_RX_BYTE_CNT_6:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_byte_cnt_6;
            REG_PORT_RX_FRAME_CNT_6:    r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_frame_cnt_6;
            REG_PORT_DIAG_STATE_6:      r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, i_port_diag_state_6};
            //REG_PORT_RX_ULTRASHORT_FRM_CNT_6: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_ultrashort_frm_cnt_6; 
            //REG_PORT_RX_OVERLENGTH_FRM_CNT_6: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_overlength_frm_cnt_6; 
            //REG_PORT_RX_CRCERR_FRM_CNT_6: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_crcerr_frm_cnt_6;     
            //REG_PORT_RX_LOOKBACK_FRM_CNT_6: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_lookback_frm_cnt_6; 
            REG_PORT_BROADFLOW_DROP_CNT_6: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_broadflow_drop_cnt_6; 
            REG_PORT_MULTIFLOW_DROP_CNT_6: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_multiflow_drop_cnt_6; 
            // �˿�8
            REG_PORT_RX_BYTE_CNT_7:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_byte_cnt_7;
            REG_PORT_RX_FRAME_CNT_7:    r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_frame_cnt_7;
            //REG_PORT_RX_FRAME_CNT_7:    r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_frame_cnt_7;
            //REG_PORT_RX_ULTRASHORT_FRM_CNT_7: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_ultrashort_frm_cnt_7; 
            //REG_PORT_RX_OVERLENGTH_FRM_CNT_7: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_overlength_frm_cnt_7; 
            //REG_PORT_RX_CRCERR_FRM_CNT_7: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_crcerr_frm_cnt_7;     
            //REG_PORT_RX_LOOKBACK_FRM_CNT_7: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_rx_lookback_frm_cnt_7; 
            //REG_PORT_BROADFLOW_DROP_CNT_7: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_broadflow_drop_cnt_7; 
            REG_PORT_MULTIFLOW_DROP_CNT_7: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_port_multiflow_drop_cnt_7; 
            // qbu_rx
            REG_QBU_RESET_0:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, r_reset_0};
            REG_RX_FRAGMENT_CNT_0:      r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_fragment_cnt_0;
            REG_RX_FRAGMENT_MISMATCH_0: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, i_rx_fragment_mismatch_0};
            REG_ERR_RX_CRC_CNT_0:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_crc_cnt_0;
            REG_ERR_RX_FRAME_CNT_0:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_frame_cnt_0;
            REG_ERR_FRAGMENT_CNT_0:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_fragment_cnt_0;
            //REG_ERR_VERIFI_CNT_0:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_verifi_cnt_0;
            REG_RX_FRAMES_CNT_0:        r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_frames_cnt_0;
            REG_FRAG_NEXT_RX_0:         r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frag_next_rx_0};
            REG_FRAME_SEQ_0:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frame_seq_0};
            
            REG_QBU_RESET_1:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, r_reset_1};
            REG_RX_FRAGMENT_CNT_1:      r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_fragment_cnt_1;
            REG_RX_FRAGMENT_MISMATCH_1: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, i_rx_fragment_mismatch_1};
            REG_ERR_RX_CRC_CNT_1:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_crc_cnt_1;
            REG_ERR_RX_FRAME_CNT_1:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_frame_cnt_1;
            REG_ERR_FRAGMENT_CNT_1:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_fragment_cnt_1;
            //REG_ERR_VERIFI_CNT_1:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_verifi_cnt_1;
            REG_RX_FRAMES_CNT_1:        r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_frames_cnt_1;
            REG_FRAG_NEXT_RX_1:         r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frag_next_rx_1};
            REG_FRAME_SEQ_1:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frame_seq_1};
            
            REG_QBU_RESET_2:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, r_reset_2};
            REG_RX_FRAGMENT_CNT_2:      r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_fragment_cnt_2;
            REG_RX_FRAGMENT_MISMATCH_2: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, i_rx_fragment_mismatch_2};
            REG_ERR_RX_CRC_CNT_2:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_crc_cnt_2;
            REG_ERR_RX_FRAME_CNT_2:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_frame_cnt_2;
            REG_ERR_FRAGMENT_CNT_2:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_fragment_cnt_2;
            //REG_ERR_VERIFI_CNT_2:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_verifi_cnt_2;
            REG_RX_FRAMES_CNT_2:        r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_frames_cnt_2;
            REG_FRAG_NEXT_RX_2:         r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frag_next_rx_2};
            REG_FRAME_SEQ_2:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frame_seq_2};
            
            REG_QBU_RESET_3:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, r_reset_3};
            REG_RX_FRAGMENT_CNT_3:      r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_fragment_cnt_3;
            REG_RX_FRAGMENT_MISMATCH_3: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, i_rx_fragment_mismatch_3};
            REG_ERR_RX_CRC_CNT_3:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_crc_cnt_3;
            REG_ERR_RX_FRAME_CNT_3:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_frame_cnt_3;
            REG_ERR_FRAGMENT_CNT_3:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_fragment_cnt_3;
            //REG_ERR_VERIFI_CNT_3:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_verifi_cnt_3;
            REG_RX_FRAMES_CNT_3:        r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_frames_cnt_3;
            REG_FRAG_NEXT_RX_3:         r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frag_next_rx_3};
            REG_FRAME_SEQ_3:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frame_seq_3};
            
            REG_QBU_RESET_4:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, r_reset_4};
            REG_RX_FRAGMENT_CNT_4:      r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_fragment_cnt_4;
            REG_RX_FRAGMENT_MISMATCH_4: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, i_rx_fragment_mismatch_4};
            REG_ERR_RX_CRC_CNT_4:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_crc_cnt_4;
            REG_ERR_RX_FRAME_CNT_4:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_frame_cnt_4;
            REG_ERR_FRAGMENT_CNT_4:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_fragment_cnt_4;
            //REG_ERR_VERIFI_CNT_4:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_verifi_cnt_4;
            REG_RX_FRAMES_CNT_4:        r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_frames_cnt_4;
            REG_FRAG_NEXT_RX_4:         r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frag_next_rx_4};
            REG_FRAME_SEQ_4:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frame_seq_4};
            
            REG_QBU_RESET_5:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, r_reset_5};
            REG_RX_FRAGMENT_CNT_5:      r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_fragment_cnt_5;
            REG_RX_FRAGMENT_MISMATCH_5: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, i_rx_fragment_mismatch_5};
            REG_ERR_RX_CRC_CNT_5:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_crc_cnt_5;
            REG_ERR_RX_FRAME_CNT_5:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_frame_cnt_5;
            REG_ERR_FRAGMENT_CNT_5:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_fragment_cnt_5;
            //REG_ERR_VERIFI_CNT_5:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_verifi_cnt_5;
            REG_RX_FRAMES_CNT_5:        r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_frames_cnt_5;
            REG_FRAG_NEXT_RX_5:         r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frag_next_rx_5};
            REG_FRAME_SEQ_5:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frame_seq_5};
            
            REG_QBU_RESET_6:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, r_reset_6};
            REG_RX_FRAGMENT_CNT_6:      r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_fragment_cnt_6;
            REG_RX_FRAGMENT_MISMATCH_6: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, i_rx_fragment_mismatch_6};
            REG_ERR_RX_CRC_CNT_6:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_crc_cnt_6;
            REG_ERR_RX_FRAME_CNT_6:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_frame_cnt_6;
            REG_ERR_FRAGMENT_CNT_6:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_fragment_cnt_6;
            //REG_ERR_VERIFI_CNT_6:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_verifi_cnt_6;
            REG_RX_FRAMES_CNT_6:        r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_frames_cnt_6;
            REG_FRAG_NEXT_RX_6:         r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frag_next_rx_6};
            REG_FRAME_SEQ_6:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frame_seq_6};
            
            REG_QBU_RESET_7:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, r_reset_7};
            REG_RX_FRAGMENT_CNT_7:      r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_fragment_cnt_7;
            REG_RX_FRAGMENT_MISMATCH_7: r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {15'd0, i_rx_fragment_mismatch_7};
            REG_ERR_RX_CRC_CNT_7:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_crc_cnt_7;
            REG_ERR_RX_FRAME_CNT_7:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_rx_frame_cnt_7;
            REG_ERR_FRAGMENT_CNT_7:     r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_fragment_cnt_7;
            //REG_ERR_VERIFI_CNT_7:       r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_err_verifi_cnt_7;
            REG_RX_FRAMES_CNT_7:        r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | i_rx_frames_cnt_7;
            REG_FRAG_NEXT_RX_7:         r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frag_next_rx_7};
            REG_FRAME_SEQ_7:            r_reg_bus_rdata <= {{REG_DATA_BUS_WIDTH{1'b0}}} | {8'd0, i_frame_seq_7};
            
            default: begin
                r_reg_bus_rdata <= {REG_DATA_BUS_WIDTH{1'b0}};
            end
        endcase
    end else begin
        r_reg_bus_rdata <= {REG_DATA_BUS_WIDTH{1'b0}};
    end
end

// �Ĵ�����������Ч��־
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_reg_bus_rdata_vld <= 1'b0;
    end else begin
        r_reg_bus_rdata_vld <= r_reg_bus_re;
    end
end

assign o_switch_reg_bus_rd_dout  = r_reg_bus_rdata;
assign o_switch_reg_bus_rd_dout_v= r_reg_bus_rdata_vld;


endmodule