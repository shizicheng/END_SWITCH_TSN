`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date: 2025/08/03 15:33:17
// Design Name: 
// Module Name: qbu_tx_timestamp
//////////////////////////////////////////////////////////////////////////////////

module qbu_tx_timestamp#(
    parameter                               DWIDTH          = 'd8                                   
)(
    input       wire                        i_clk                       ,
    input       wire                        i_rst                       ,

    input       wire    [DWIDTH - 1:0]      i_mac_axis_data             ,          
    input       wire                        i_mac_axis_valid            ,              

    output      wire                        o_mac_time_irq              , // ��ʱ����ж��ź�
    output      wire    [7:0]               o_mac_frame_seq             , // ֡���к�
    output      wire    [7:0]               o_timestamp_addr              // ��ʱ����洢�� RAM ��ַ
);

    //==========================================================================
    // ��������
    //==========================================================================
    localparam                              PTP_ETHERTYPE   = 16'h88F7  ; // PTP Э������
    localparam                              BYTE_CNT_WIDTH  = 'd8       ; // �ֽڼ�����λ��

    //==========================================================================
    // �����źżĴ��� (ri_ ��ͷ)
    //==========================================================================
    reg         [DWIDTH - 1:0]              ri_mac_axis_data            ;
    reg                                     ri_mac_axis_valid           ;

    //==========================================================================
    // �ڲ��߼��ź�
    //==========================================================================
    wire                                    w_data_valid                ; // ������Ч�ź�
    wire                                    w_frame_start               ; // ֡��ʼ�ź�
    wire                                    w_ptp_ethertype_match       ; // PTP ��̫������ƥ��
    wire                                    w_ptp_trigger               ; // PTP ʱ�����������
    
    //==========================================================================
    // �ڲ��Ĵ���
    //==========================================================================
    reg         [BYTE_CNT_WIDTH-1:0]        r_byte_counter              ; // �ֽڼ�����
    reg         [15:0]                      r_ethertype_buffer          ; // ��̫�����ͻ���
    reg                                     r_ptp_frame_flag            ; // PTP ���ı�־
    reg         [7:0]                       r_ptp_message_type          ; // PTP ��Ϣ���ͻ���
    reg                                     r_data_valid_d1             ; // ������Ч�ź��ӳ�һ��

    //==========================================================================
    // ����źżĴ��� (ro_ ��ͷ)
    //==========================================================================
    reg                                     ro_mac_time_irq             ;
    reg         [7:0]                       ro_mac_frame_seq            ;
    reg         [7:0]                       ro_timestamp_addr           ;

    //==========================================================================
    // �����źżĴ�
    //==========================================================================
    always @(posedge i_clk or posedge i_rst) begin
        if (i_rst) begin
            ri_mac_axis_data            <= {DWIDTH{1'b0}} ;
            ri_mac_axis_valid           <= 1'b0    ;
        end else begin
            ri_mac_axis_data            <= i_mac_axis_data ;
            ri_mac_axis_valid           <= i_mac_axis_valid;
        end
    end

    //==========================================================================
    // ����߼�
    //==========================================================================
    // ������Ч�ź�
    assign w_data_valid = ri_mac_axis_valid;
    
    // ֡��ʼ��⣺��Ч������ǰһ����Ч
    assign w_frame_start = w_data_valid && (~r_data_valid_d1);
    
    // PTP ��̫������ƥ��
    assign w_ptp_ethertype_match = (r_ethertype_buffer == PTP_ETHERTYPE);
    
    // PTP ʱ�������������PTP ��������Ϣ����[3:0]Ϊ 0x0, 0x2, 0x3
    assign w_ptp_trigger = r_ptp_frame_flag && (r_byte_counter == 8'd11) && w_data_valid &&
                          ((ri_mac_axis_data[3:0] == 4'h0) || 
                           (ri_mac_axis_data[3:0] == 4'h2) || 
                           (ri_mac_axis_data[3:0] == 4'h3));

    //==========================================================================
    // ʱ���߼�
    //==========================================================================
    // ������Ч�ź��ӳ�
    always @(posedge i_clk or posedge i_rst) begin
        if (i_rst) begin
            r_data_valid_d1 <= 1'b0;
        end else begin
            r_data_valid_d1 <= w_data_valid;
        end
    end

    // �ֽڼ�������ÿ֡��0��ʼ����
    always @(posedge i_clk or posedge i_rst) begin
        if (i_rst) begin
            r_byte_counter <= 8'd0;
        end else if (w_frame_start) begin
            r_byte_counter <= 8'd1;
        end else if (w_data_valid) begin
            r_byte_counter <= r_byte_counter + 1'b1;
        end
    end

    // ��̫�����ͻ��棺�����9��10�ֽ�
    always @(posedge i_clk or posedge i_rst) begin
        if (i_rst) begin
            r_ethertype_buffer <= 16'd0;
        end else if (w_data_valid) begin
            if (r_byte_counter == 8'd9) begin
                r_ethertype_buffer[15:8] <= ri_mac_axis_data;
            end else if (r_byte_counter == 8'd10) begin
                r_ethertype_buffer[7:0] <= ri_mac_axis_data;
            end
        end
    end

    // PTP ���ı�־����⵽PTP��̫�����ͺ���λ��֡����������
    always @(posedge i_clk or posedge i_rst) begin
        if (i_rst) begin
            r_ptp_frame_flag <= 1'b0;
        end else if (w_frame_start) begin
            r_ptp_frame_flag <= 1'b0;
        end else if ((r_byte_counter == 8'd10) && w_data_valid && w_ptp_ethertype_match) begin
            r_ptp_frame_flag <= 1'b1;
        end
    end

    // PTP ��Ϣ���ͻ��棺�����11�ֽ�
    always @(posedge i_clk or posedge i_rst) begin
        if (i_rst) begin
            r_ptp_message_type <= 8'd0;
        end else if (w_data_valid && (r_byte_counter == 8'd11)) begin
            r_ptp_message_type <= ri_mac_axis_data;
        end
    end

    // ֡���кż�������ÿ���յ�һ����Ч����֡���кż�1
    always @(posedge i_clk or posedge i_rst) begin
        if (i_rst) begin
            ro_mac_frame_seq <= 8'd0;
        end else if (w_data_valid) begin
            ro_mac_frame_seq <= ro_mac_frame_seq + 1'b1;
        end
    end

    // ʱ����ж��źţ����� PTP ��������ʱ����
    always @(posedge i_clk or posedge i_rst) begin
        if (i_rst) begin
            ro_mac_time_irq <= 1'b0;
        end else begin
            ro_mac_time_irq <= w_ptp_trigger;
        end
    end

    // ʱ�����ַ��������ÿ�β���ʱ����ж�ʱ��ַ��1
    always @(posedge i_clk or posedge i_rst) begin
        if (i_rst) begin
            ro_timestamp_addr <= 8'd0;
        end else if (w_ptp_trigger) begin
            ro_timestamp_addr <= ro_timestamp_addr + 1'b1;
        end
    end

    //==========================================================================
    // ����źŸ�ֵ
    //==========================================================================
    assign o_mac_time_irq       = ro_mac_time_irq      ;
    assign o_mac_frame_seq      = ro_mac_frame_seq     ;
    assign o_timestamp_addr     = ro_timestamp_addr    ;

endmodule
