`include "synth_cmd_define.vh"

module  Scheduling_top #(
    parameter                                                   PORT_FIFO_PRI_NUM       =      8    ,  // ֧�ֶ˿����ȼ� FIFO ������
    parameter                                                   REG_ADDR_BUS_WIDTH      =      8    ,
    parameter                                                   REG_DATA_BUS_WIDTH      =      16     
)(
    input               wire                                    i_clk                            , // 250MHz
    input               wire                                    i_rst                            ,
    /*----------- �Ĵ������ýӿ� ------------*/
    // �Ĵ��������ź�                     
    //input               wire                                    i_refresh_list_pulse             , // ˢ�¼Ĵ����б�״̬�Ĵ����Ϳ��ƼĴ�����
    //input               wire                                    i_switch_err_cnt_clr             , // ˢ�´��������
    //input               wire                                    i_switch_err_cnt_stat            , // ˢ�´���״̬�Ĵ���
    // �Ĵ���д���ƽӿ�     
    //input               wire                                    i_Sch_reg_bus_we                 , // �Ĵ���дʹ��
    //input               wire   [REG_ADDR_BUS_WIDTH-1:0]         i_Sch_reg_bus_we_addr            , // �Ĵ���д��ַ
    //input               wire   [REG_DATA_BUS_WIDTH-1:0]         i_Sch_reg_bus_we_din             , // �Ĵ���д����
    //input               wire                                    i_Sch_reg_bus_we_din_v           , // �Ĵ���д����ʹ��
    // �Ĵ��������ƽӿ�     
    //input               wire                                    i_Sch_reg_bus_rd                 , // �Ĵ�����ʹ��
    //input               wire   [REG_ADDR_BUS_WIDTH-1:0]         i_Sch_reg_bus_rd_addr            , // �Ĵ�������ַ
    //output              wire   [REG_DATA_BUS_WIDTH-1:0]         o_Sch_reg_bus_we_dout            , // �����Ĵ�������
    //output              wire                                    o_Sch_reg_bus_we_dout_v          , // ��������Чʹ��
    /*------------------------------------ Schedule�Ĵ��� ----------------------------------------*/
    input               wire   [7:0]                            i_idleSlope_q0             			,
    input               wire   [7:0]                            i_idleSlope_q1             			,
    input               wire   [7:0]                            i_idleSlope_q2             			,
    input               wire   [7:0]                            i_idleSlope_q3             			,
    input               wire   [7:0]                            i_idleSlope_q4             			,
    input               wire   [7:0]                            i_idleSlope_q5             			,
    input               wire   [7:0]                            i_idleSlope_q6             			,
    input               wire   [7:0]                            i_idleSlope_q7             			,
	input   			wire   [7:0]                            i_sendslope_q0             			,
    input               wire   [7:0]                            i_sendslope_q1             			,
    input               wire   [7:0]                            i_sendslope_q2             			,
    input               wire   [7:0]                            i_sendslope_q3             			,
    input               wire   [7:0]                            i_sendslope_q4             			,
    input               wire   [7:0]                            i_sendslope_q5             			,
    input               wire   [7:0]                            i_sendslope_q6             			,
    input               wire   [7:0]                            i_sendslope_q7             			,
	input   			wire                                    i_qav_en                 			,
	input   			wire   [15:0]                           i_lothreshold_q0             	    ,
    input               wire   [15:0]                           i_lothreshold_q1             		,
    input               wire   [15:0]                           i_lothreshold_q2             		,
    input               wire   [15:0]                           i_lothreshold_q3           			,
    input               wire   [15:0]                           i_lothreshold_q4           			,
    input               wire   [15:0]                           i_lothreshold_q5           			,
    input               wire   [15:0]                           i_lothreshold_q6           			,
    input               wire   [15:0]                           i_lothreshold_q7           			,
    input               wire   [15:0]                           i_hithreshold_q0           			,
    input               wire   [15:0]                           i_hithreshold_q1           			,
    input               wire   [15:0]                           i_hithreshold_q2           			,
    input               wire   [15:0]                           i_hithreshold_q3           			,
    input               wire   [15:0]                           i_hithreshold_q4           			,
    input               wire   [15:0]                           i_hithreshold_q5           			,
    input               wire   [15:0]                           i_hithreshold_q6           			,
    input               wire   [15:0]                           i_hithreshold_q7           			,
    
	input   			wire                                    i_config_vld             			,


    input               wire   [79:0]                           i_current_time                      ,
	input   			wire   [79:0]                           i_Base_time              			, 
	input   			wire                                    i_ConfigChange           			,
	input   			wire   [PORT_FIFO_PRI_NUM-1:0]          i_ControlList            			,     
	input   			wire   [7:0]                            i_ControlList_len        			,    
	input   			wire                                    i_ControlList_vld        			,     
	input   			wire   [15:0]                           i_cycle_time             			,    
	input   			wire   [79:0]                           i_cycle_time_extension   			, 
	input   			wire                                    i_qbv_en                 			,       
			  		  
	input   			wire   [3:0]                            i_qos_sch                           ,
	input   			wire	                                i_qos_en                            ,   

    /*------------------------------ ��CROSSBAR����ƽ�潻���ĵ�����Ϣ ------------------------------*/
    // ������ˮ�ߵ�����Ϣ����
    input               wire  [PORT_FIFO_PRI_NUM-1:0]           i_fifoc_empty                       , // ʵʱ���ö˿ڶ�Ӧ CROSSBAR ����ƽ�����ȼ� FIFO ��Ϣ 
    output              wire  [PORT_FIFO_PRI_NUM-1:0]           o_scheduing_rst                     , // �ö˿ڵ�����ˮ�߲����ĵ��Ƚ��
    output              wire                                    o_scheduing_rst_vld                 , // �ö˿ڵ�����ˮ�߲����ĵ��Ƚ����Чλ
    // QBU ģ�鷵�ص��ź�
    input               wire                                    i_mac_tx_axis_valid                 , // ���ڹ���ÿ�����ȼ����е�����ֵ
    input               wire                                    i_mac_tx_axis_last                  ,  // ������ last �źţ�����ʹ�ܵ�����ˮ�߼���  
    input               wire  [15:0]                            i_mac_tx_axis_user
);

/*------------ wire -----------*/
wire   [PORT_FIFO_PRI_NUM-1:0]          w_queque                 ;
wire                                    w_queque_vld             ;
 
wire   [PORT_FIFO_PRI_NUM-1:0]          w_ControlList_state      ;
wire                                    w_ControlList_state_vld  ;
 
wire   [PORT_FIFO_PRI_NUM-1:0]          w_qos_scheduing_res      ;
wire                                    w_qos_scheduing_rst_vld  ;
/*
wire   [7:0]                            w_idleSlope              ;
wire   [7:0]                            w_sendslope              ;
wire                                    w_qav_en                 ;
wire   [15:0]                           w_threshold              ;
wire                                    w_config_vld             ;

wire   [79:0]                           w_Base_time              ; 
wire                                    w_ConfigChange           ;
wire   [PORT_FIFO_PRI_NUM:0]            w_ControlList            ;     
wire   [7:0]                            w_ControlList_len        ;    
wire                                    w_ControlList_vld        ;     
wire   [15:0]                           w_cycle_time             ;    
wire   [79:0]                           w_cycle_time_extension   ; 
wire                                    w_qbv_en                 ;       
 
wire   [3:0]                            w_qos_sch                ;
wire                                    w_qos_en                 ;                         
*/
tsn_qav_mng #(
    .PORT_FIFO_PRI_NUM       ( PORT_FIFO_PRI_NUM       )      // ֧�ֶ˿����ȼ� FIFO ������
) tsn_qav_mng_inst ( 
    .i_clk                   ( i_clk                   ) , // 250MHz
    .i_rst                   ( i_rst                   ) ,
    /*------------------------------ �Ĵ������ýӿ� ----------------------------*/
    .i_idleSlope_q0           ( i_idleSlope_q0            ) ,
    .i_idleSlope_q1           ( i_idleSlope_q1            ) ,
    .i_idleSlope_q2           ( i_idleSlope_q2            ) ,
    .i_idleSlope_q3           ( i_idleSlope_q3            ) ,
    .i_idleSlope_q4           ( i_idleSlope_q4            ) ,
    .i_idleSlope_q5           ( i_idleSlope_q5            ) ,
    .i_idleSlope_q6           ( i_idleSlope_q6            ) ,
    .i_idleSlope_q7           ( i_idleSlope_q7            ) ,
    .i_sendslope_q0           ( i_sendslope_q0          ) ,
    .i_sendslope_q1           ( i_sendslope_q1          ) ,
    .i_sendslope_q2           ( i_sendslope_q2          ) ,
    .i_sendslope_q3           ( i_sendslope_q3          ) ,
    .i_sendslope_q4           ( i_sendslope_q4          ) ,
    .i_sendslope_q5           ( i_sendslope_q5          ) ,
    .i_sendslope_q6           ( i_sendslope_q6          ) ,
    .i_sendslope_q7           ( i_sendslope_q7          ) ,
    .i_hithreshold_q0           ( i_hithreshold_q0          ) ,
    .i_hithreshold_q1           ( i_hithreshold_q1          ) ,
    .i_hithreshold_q2           ( i_hithreshold_q2          ) ,
    .i_hithreshold_q3           ( i_hithreshold_q3          ) ,
    .i_hithreshold_q4           ( i_hithreshold_q4          ) ,
    .i_hithreshold_q5           ( i_hithreshold_q5          ) ,
    .i_hithreshold_q6           ( i_hithreshold_q6          ) ,
    .i_hithreshold_q7           ( i_hithreshold_q7          ) ,
    .i_lothreshold_q0           ( i_lothreshold_q0          ) ,
    .i_lothreshold_q1           ( i_lothreshold_q1          ) ,
    .i_lothreshold_q2           ( i_lothreshold_q2          ) ,
    .i_lothreshold_q3           ( i_lothreshold_q3          ) ,
    .i_lothreshold_q4           ( i_lothreshold_q4          ) ,
    .i_lothreshold_q5           ( i_lothreshold_q5          ) ,
    .i_lothreshold_q6           ( i_lothreshold_q6          ) ,
    .i_lothreshold_q7           ( i_lothreshold_q7          ) ,
    
    .i_config_vld            ( i_config_vld            ) ,
    .i_qav_en                ( i_qav_en                ) ,
    /*------------------------------ ������Ϣ���� ------------------------------*/
    .i_fifoc_empty           ( i_fifoc_empty           ) , // ʵʱ���ö˿ڶ�Ӧ CROSSBAR ����ƽ�����ȼ� FIFO ��Ϣ
    .i_scheduing_rst         ( w_qos_scheduing_res     ) , // �ö˿ڵ�����ˮ�߲����ĵ��Ƚ��
    .i_scheduing_rst_vld     ( w_qos_scheduing_rst_vld ) , // �ö˿ڵ�����ˮ�߲����ĵ��Ƚ����Чλ
    .i_mac_tx_axis_valid     ( i_mac_tx_axis_valid     ) , // ���ڹ���ÿ�����ȼ����е�����ֵ
    .i_mac_tx_axis_last      ( i_mac_tx_axis_last      ) , // 
    .i_mac_tx_axis_user      ( i_mac_tx_axis_user      ) ,
    /*---------------- ������ֵ���������������ȼ�������Ϣ��� ------------------*/
    .o_queue                ( w_queque                ) , // �����������ֵ�Ķ��н������
    .o_queue_vld            ( w_queque_vld            ) 
);

tsn_qbv_mng #(
    .PORT_FIFO_PRI_NUM       (PORT_FIFO_PRI_NUM       )      // ֧�ֶ˿����ȼ� FIFO ������
) tsn_qbv_mng_inst ( 
    .i_clk                   ( i_clk                  ) , // 250MHz
    .i_rst                   ( i_rst                  ) ,
    /*---------------------------------------- �Ĵ������ýӿ� --------------------------------------*/
    .i_current_time          ( i_current_time         ) ,
    .i_Base_time             ( i_Base_time            ) ,
    .i_Base_time_vld         ( 1'b0                   ),
    .i_ConfigChange          ( i_ConfigChange         ) ,
    .i_ControlList           ( i_ControlList          ) ,   
    .i_ControlList_len       ( i_ControlList_len      ) , 
    .i_ControlList_vld       ( i_ControlList_vld      ) ,   
    .i_cycle_time            ( i_cycle_time           ) ,      
    .i_cycle_time_extension  ( i_cycle_time_extension ) ,
    .i_qbv_en                ( i_qbv_en               ) ,  
    /*---------------------------------- Qav �����������������Ķ���������� -------------------------*/ 
    .i_queque                ( w_queque               ) , // �����������ֵ�Ķ��н������
    .i_queque_vld            ( w_queque_vld           ) ,
    /*---------------------------------- ����ſ�״̬�� QOS ����ģ�� ------------------------------*/ 
    .o_ControlList_state     ( w_ControlList_state    ) , // �ſ��б��״̬
    .o_ControlList_state_vld ( w_ControlList_state_vld) 
);

tx_qos_mng #(
    .PORT_FIFO_PRI_NUM       ( PORT_FIFO_PRI_NUM       )                       // ֧�ֶ˿����ȼ� FIFO ������
)tx_qos_mng_inst(   
    .i_clk                   ( i_clk                   ) ,   // 250MHz
    .i_rst                   ( i_rst                   ) ,
    /*---------------------------------------- �Ĵ������ýӿ� -------------------------------------------*/
    .i_qos_sch               ( i_qos_sch               ) ,
    .i_qos_en                ( i_qos_en                ) ,
    /*---------------------------- ���ݵ����㷨�����Ҫ�������ȼ����� --------------------------------*/ 
    .i_ControlList_state     ( w_ControlList_state     ) ,  // �ſ��б��״̬
    .i_qos_req               ( w_ControlList_state_vld ) ,
    .o_qos_scheduing_res     ( w_qos_scheduing_res     ) ,
    .o_qos_scheduing_rst_vld ( w_qos_scheduing_rst_vld )                 
);

assign o_scheduing_rst     = w_qos_scheduing_res;
assign o_scheduing_rst_vld = w_qos_scheduing_rst_vld;

/*
Schduling_regs #(
    .PORT_FIFO_PRI_NUM       ( PORT_FIFO_PRI_NUM  )  ,  // ֧�ֶ˿����ȼ� FIFO ������
    .REG_ADDR_BUS_WIDTH      ( REG_ADDR_BUS_WIDTH )  ,
    .REG_DATA_BUS_WIDTH      ( REG_DATA_BUS_WIDTH )    
) Schduling_regs_inst (
    .i_clk                   ( i_clk                   )        ,
    .i_rst                   ( i_rst                   )        ,
    // �Ĵ������ýӿ�
    // �Ĵ��������ź�                     
    .i_refresh_list_pulse    ( i_refresh_list_pulse    )        , // ˢ�¼Ĵ����б�״̬�Ĵ����Ϳ��ƼĴ�����
    .i_switch_err_cnt_clr    ( i_switch_err_cnt_clr    )        , // ˢ�´��������
    .i_switch_err_cnt_stat   ( i_switch_err_cnt_stat   )        , // ˢ�´���״̬�Ĵ���
    // �Ĵ���д���ƽӿ�     
    .i_Sch_reg_bus_we        ( i_Sch_reg_bus_we        )        , // �Ĵ���дʹ��
    .i_Sch_reg_bus_we_addr   ( i_Sch_reg_bus_we_addr   )        , // �Ĵ���д��ַ
    .i_Sch_reg_bus_we_din    ( i_Sch_reg_bus_we_din    )        , // �Ĵ���д����
    .i_Sch_reg_bus_we_din_v  ( i_Sch_reg_bus_we_din_v  )        , // �Ĵ���д����ʹ��
    // �Ĵ��������ƽӿ�     
    .i_Sch_reg_bus_rd        ( i_Sch_reg_bus_rd        )         , // �Ĵ�����ʹ��
    .i_Sch_reg_bus_rd_addr   ( i_Sch_reg_bus_rd_addr   )         , // �Ĵ�������ַ
    .o_Sch_reg_bus_we_dout   ( o_Sch_reg_bus_we_dout   )         , // �����Ĵ�������
    .o_Sch_reg_bus_we_dout_v ( o_Sch_reg_bus_we_dout_v )         , // ��������Чʹ��
    // IP�����������Ϣ
    // qav
    .o_idleSlope             ( w_idleSlope            )         ,
    .o_sendslope             ( w_sendslope            )         ,
    .o_qav_en                ( w_qav_en               )         ,
    .o_threshold             ( w_threshold            )         ,  
    .o_av_config_vld         ( w_config_vld           )         ,
    // qbv
    .o_Base_time             ( w_Base_time            )         ,
    .o_ConfigChange          ( w_ConfigChange         )         ,
    .o_ControlList           ( w_ControlList          )         ,   
    .o_ControlList_len       ( w_ControlList_len      )         ,  
    .o_ControlList_vld       ( w_ControlList_vld      )         ,
    .o_cycle_time            ( w_cycle_time           )         ,      
    .o_cycle_time_extension  ( w_cycle_time_extension )         ,
    .o_qbv_en                ( w_qbv_en               )         ,       
    // qos 
    .o_qos_sch               ( w_qos_sch              )         ,
    .o_qos_en                ( w_qos_en               )                                  
);
*/
endmodule