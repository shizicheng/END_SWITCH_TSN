module rx_port_mng#(
    parameter                                                   PORT_NUM                =      4        ,  // �������Ķ˿���
    parameter                                                   PORT_MNG_DATA_WIDTH     =      8        ,  // Mac_port_mng ����λ��
    parameter                                                   HASH_DATA_WIDTH         =      15       ,  // ��ϣ�����ֵ��λ�� 
    parameter                                                   REG_ADDR_BUS_WIDTH      =      8        ,  // ���� MAC ������üĴ�����ַλ��
    parameter                                                   REG_DATA_BUS_WIDTH      =      16       ,  // ���� MAC ������üĴ�������λ��
    parameter                                                   METADATA_WIDTH          =      94       ,  // ��Ϣ��λ��
    parameter                                                   LOOK_UP_DATA_WIDTH      =      144      ,  // ����ͷ��Ϣ MAC + VLAN + Eth_type
    parameter                                                   CAM_NUM                 =      256      ,
    parameter                                                   CROSS_DATA_WIDTH        =     PORT_MNG_DATA_WIDTH, // �ۺ��������
    parameter                                                   PORT_FIFO_PRI_NUM       =      8        ,  // ���ȼ�FIFO����
    parameter   [31:0]                                          PORT_INDEX              =      32'd0       // �˿���������
)(
    input               wire                                    i_clk                              ,   // 250MHz
    input               wire                                    i_rst                              ,
    
    // �Ĵ��������ź�
    //input               wire                                    i_refresh_list_pulse                , // ˢ�¼Ĵ����б�״̬�Ĵ����Ϳ��ƼĴ�����
    //input               wire                                    i_switch_err_cnt_clr                , // ˢ�´��������
    //input               wire                                    i_switch_err_cnt_stat               , // ˢ�´���״̬�Ĵ���
    // �Ĵ���д���ƽӿ�
    //input               wire                                    i_switch_reg_bus_we                , // �Ĵ���дʹ��
    //input               wire   [REG_ADDR_BUS_WIDTH-1:0]         i_switch_reg_bus_we_addr           , // �Ĵ���д��ַ
    //input               wire   [REG_DATA_BUS_WIDTH-1:0]         i_switch_reg_bus_we_din            , // �Ĵ���д����
    //input               wire                                    i_switch_reg_bus_we_din_v          , // �Ĵ���д����ʹ��
    // �Ĵ��������ƽӿ�
    //input               wire                                    i_switch_reg_bus_rd                , // �Ĵ�����ʹ��
    //input               wire   [REG_ADDR_BUS_WIDTH-1:0]         i_switch_reg_bus_rd_addr           , // �Ĵ�������ַ
    //output              wire   [REG_DATA_BUS_WIDTH-1:0]         o_switch_reg_bus_we_dout           , // �����Ĵ�������
    //output              wire                                    o_switch_reg_bus_we_dout_v         , // ��������Чʹ��
    
    /*---------------------------------------- ����� MAC ������ -------------------------------------------*/
    input               wire                                    i_mac_port_link                    , // �˿ڵ�����״̬
    input               wire   [1:0]                            i_mac_port_speed                   , // �˿�������Ϣ��00-10M��01-100M��10-1000M��10-10G
    input               wire                                    i_mac_port_filter_preamble_v       , // �˿��Ƿ����ǰ������Ϣ
    input               wire   [PORT_MNG_DATA_WIDTH-1:0]        i_mac_axi_data                     , // �˿�������
    input               wire   [(PORT_MNG_DATA_WIDTH/8)-1:0]    i_mac_axi_data_keep                , // �˿����������룬��Ч�ֽ�ָʾ
    input               wire                                    i_mac_axi_data_valid               , // �˿�������Ч
    output              wire                                    o_mac_axi_data_ready               , // �˿����ݾ����ź�,��ʾ��ǰģ��׼���ý�������
    input               wire                                    i_mac_axi_data_last                , // ������������ʶ
    //ʱ����ź�
	output              wire                                    o_mac_time_irq                     , // ��ʱ����ж��ź�
    output              wire   [7:0]                            o_mac_frame_seq                    , // ֡���к�
    output              wire   [6:0]                            o_timestamp_addr                   ,  // ��ʱ����洢�� RAM ��ַ
    /*---------------------------------------- ����Ĺ�ϣֵ -------------------------------------------*/ 
    output              wire   [11:0]                           o_vlan_id                          ,
    output              wire   [HASH_DATA_WIDTH - 1 : 0]        o_dmac_hash_key                    , // Ŀ�� mac �Ĺ�ϣֵ
    output              wire   [47 : 0]                         o_dmac                             , // Ŀ�� mac ��ֵ
    output              wire                                    o_dmac_vld                         , // dmac_vld
    output              wire   [HASH_DATA_WIDTH - 1 : 0]        o_smac_hash_key                    , // Դ mac ��ֵ��Ч��ʶ
    output              wire   [47 : 0]                         o_smac                             , // Դ mac ��ֵ
    output              wire                                    o_smac_vld                         , // smac_vld
    /*---------------------------------------- ���ҵ�ת���˿ں� ---------------------------------------*/
    input               wire   [PORT_NUM-1:0]                   i_swlist_tx_port                   , // �������Ͷ˿���Ϣ
    input               wire                                    i_swlist_vld                       , // ���Ͷ˿��ź���Ч�ź� 
    input               wire   [1:0]                            i_swlist_port_broadcast            , // 01:�鲥 10���㲥 11:����
    // ���潻���߼�
    output             wire                                     o_rtag_flag                        , // �Ƿ�Я��rtag��ǩ,��CBҵ��֡,��Ҫ�ȹ�CBģ������Ƿ�����,������crossbar
    output             wire   [15:0]                            o_rtag_squence                     , // rtag_squencenum
    output             wire   [7:0]                             o_stream_handle                    , // ACL��ʶ��,��������ÿ��������ά���Լ���

    input              wire                                     i_pass_en                          , // �жϽ�������Խ��ո�֡
    input              wire                                     i_discard_en                       , // �жϽ�������Զ�����֡
    input              wire                                     i_judge_finish                     , // �жϽ������ʾ���α��ĵ��ж����  

    output             wire                                     o_tx_req                           ,
    input              wire                                     i_mac_tx0_ack                      , // ��Ӧʹ���ź�
    input              wire   [PORT_FIFO_PRI_NUM-1:0]           i_mac_tx0_ack_rst                  , // �˿ڵ����ȼ��������
    input              wire                                     i_mac_tx1_ack                      , // ��Ӧʹ���ź�
    input              wire   [PORT_FIFO_PRI_NUM-1:0]           i_mac_tx1_ack_rst                  , // �˿ڵ����ȼ��������  
    input              wire                                     i_mac_tx2_ack                      , // ��Ӧʹ���ź�
    input              wire   [PORT_FIFO_PRI_NUM-1:0]           i_mac_tx2_ack_rst                  , // �˿ڵ����ȼ��������
    input              wire                                     i_mac_tx3_ack                      , // ��Ӧʹ���ź�
    input              wire   [PORT_FIFO_PRI_NUM-1:0]           i_mac_tx3_ack_rst                  , // �˿ڵ����ȼ��������
    input              wire                                     i_mac_tx4_ack                      , // ��Ӧʹ���ź�
    input              wire   [PORT_FIFO_PRI_NUM-1:0]           i_mac_tx4_ack_rst                  , // �˿ڵ����ȼ��������
    input              wire                                     i_mac_tx5_ack                      , // ��Ӧʹ���ź�
    input              wire   [PORT_FIFO_PRI_NUM-1:0]           i_mac_tx5_ack_rst                  , // �˿ڵ����ȼ��������
    input              wire                                     i_mac_tx6_ack                      , // ��Ӧʹ���ź�
    input              wire   [PORT_FIFO_PRI_NUM-1:0]           i_mac_tx6_ack_rst                  , // �˿ڵ����ȼ��������
    input              wire                                     i_mac_tx7_ack                      , // ��Ӧʹ���ź�
    input              wire   [PORT_FIFO_PRI_NUM-1:0]           i_mac_tx7_ack_rst                  , // �˿ڵ����ȼ��������


    /*---------------------------------------- �� PORT ��������� -------------------------------------------*/
    output              wire                                    o_mac_cross_port_link              , // �˿ڵ�����״̬
    output              wire   [1:0]                            o_mac_cross_port_speed             , // �˿�������Ϣ��00-10M��01-100M��10-1000M��10-10G 
    output              wire   [CROSS_DATA_WIDTH-1:0]           o_mac_cross_port_axi_data          , // �˿������������λ��ʾcrcerr
    output              wire   [15:0]                           o_mac_cross_port_axi_user          ,
    output              wire   [(CROSS_DATA_WIDTH/8)-1:0]       o_mac_cross_axi_data_keep          , // �˿����������룬��Ч�ֽ�ָʾ
    output              wire                                    o_mac_cross_axi_data_valid         , // �˿�������Ч
    input               wire                                    i_mac_cross_axi_data_ready         , // �������߾ۺϼܹ���ѹ��ˮ���ź�
    output              wire                                    o_mac_cross_axi_data_last          , // ������������ʶ
    /*---------------------------------------- �� PORT �ۺ���Ϣ�� -------------------------------------------*/
    output             wire   [METADATA_WIDTH-1:0]              o_cross_metadata                   , // ���� metadata ����
    output             wire                                     o_cross_metadata_valid             , // ���� metadata ������Ч�ź�
    output             wire                                     o_cross_metadata_last              , // ��Ϣ��������ʶ
    input              wire                                     i_cross_metadata_ready             , // ����ģ�鷴ѹ��ˮ�� 
    /*---------------------------------------- �� PORT �ؼ�֡��������� -------------------------------------------*/ 
    output              wire   [CROSS_DATA_WIDTH-1:0]           o_emac_port_axi_data               , // �˿������������λ��ʾcrcerr
    output              wire   [15:0]                           o_emac_port_axi_user               ,
    output              wire   [(CROSS_DATA_WIDTH/8)-1:0]       o_emac_axi_data_keep               , // �˿����������룬��Ч�ֽ�ָʾ
    output              wire                                    o_emac_axi_data_valid              , // �˿�������Ч
    input               wire                                    i_emac_axi_data_ready              , // �������߾ۺϼܹ���ѹ��ˮ���ź�
    output              wire                                    o_emac_axi_data_last               , // ������������ʶ
    /*---------------------------------------- �� PORT �ۺ���Ϣ�� -------------------------------------------*/
    output              wire   [METADATA_WIDTH-1:0]             o_emac_metadata                    , // ���� metadata ����
    output              wire                                    o_emac_metadata_valid              , // ���� metadata ������Ч�ź�
    output              wire                                    o_emac_metadata_last               , // ��Ϣ��������ʶ
    input               wire                                    i_emac_metadata_ready              , // ����ģ�鷴ѹ��ˮ�� 
/*
        metadata �������
            
            [80:65] : CBЭ�� R-TAG�ֶ� ok
            [64:63](2bit) : port_speed ok
            [62:60](3bit) : vlan_pri ok
            [59:52](8bit) : tx_prot ok 
            [51:44](8bit) : acl_frmtype ok
            [43:28](16bit): acl_fetchinfo ok
            [27](1bit) : frm_vlan_flag ok
            [26:19](8bit) : ����˿ڣ�bitmap��ʾ ok
            [18:15](4bit) : ����
            [14:13](2bit) : ��ʶ��ƥ�䣬[0]:1��ʾCBҵ��֡��[0]:0��ʾ��CBҵ��֡  [1]��1 �� rtag ��ǩ [1]��0 �� rtag ��ǩ ok 
            [12](1bit) : ����λ ok
            [11](1bit) : �Ƿ�Ϊ�ؼ�֡(Qbu)  ok
            [10:4](7bit) ��time_stamp_addr������ʱ����ĵ�ַ��Ϣ  ok
            [3:0](3bit): ����
    */
    //qbu��֤�ź�
    output             wire                                     o_qbu_verify_valid                 ,
    output             wire                                     o_qbu_response_valid               ,

    /*---------------------------------------- ƽ̨�Ĵ��������� RXMAC ��صļĴ��� -------------------------------------------*/
    input              wire   [15:0]                            i_hash_ploy_regs                   , // ��ϣ����ʽ
    input              wire   [15:0]                            i_hash_init_val_regs               , // ��ϣ����ʽ��ʼֵ
    input              wire                                     i_hash_regs_vld                    ,
    input              wire                                     i_port_rxmac_down_regs             , // �˿ڽ��շ���MAC�ر�ʹ��
    input              wire                                     i_port_broadcast_drop_regs         , // �˿ڹ㲥֡����ʹ��
    input              wire                                     i_port_multicast_drop_regs         , // �˿��鲥֡����ʹ��
    input              wire                                     i_port_loopback_drop_regs          , // �˿ڻ���֡����ʹ��
    input              wire   [47:0]                            i_port_mac_regs                    , // �˿ڵ� MAC ��ַ
    input              wire                                     i_port_mac_vld_regs                , // ʹ�ܶ˿� MAC ��ַ��Ч
    input              wire   [7:0]                             i_port_mtu_regs                    , // MTU����ֵ
    input              wire   [PORT_NUM-1:0]                    i_port_mirror_frwd_regs            , // ����ת���Ĵ���������Ӧ�Ķ˿���1���򱾶˿ڽ��յ����κ�ת������֡������ת��ֵ����1�Ķ˿�
    input              wire   [15:0]                            i_port_flowctrl_cfg_regs           , // ������������
    input              wire   [4:0]                             i_port_rx_ultrashortinterval_num   , // ֡���
    // ACL �Ĵ���
    input              wire   [PORT_NUM-1:0]                    i_acl_port_sel                     , // ѡ��Ҫ���õĶ˿�
	input			   wire										i_acl_port_sel_valid			   ,
    input              wire                                     i_acl_clr_list_regs                , // ��ռĴ����б�
    output             wire                                     o_acl_list_rdy_regs                , // ���üĴ�����������
    input              wire   [4:0]                             i_acl_item_sel_regs                , // ������Ŀѡ��
// DMAC����ֵ���ã�6��16λ�ֶΣ�
    input    			wire [15:0]                      		i_cfg_acl_item_dmac_code_1            , // �˿�ACL����-д��dmacֵ[15:0]
    input    			wire                             		i_cfg_acl_item_dmac_code_1_valid      , // д����Ч�ź�
					
    input    			wire [15:0]                      		i_cfg_acl_item_dmac_code_2            , // �˿�ACL����-д��dmacֵ[31:16]
    input    			wire                             		i_cfg_acl_item_dmac_code_2_valid      , // д����Ч�ź�
					
    input    			wire [15:0]                      		i_cfg_acl_item_dmac_code_3            , // �˿�ACL����-д��dmacֵ[47:32]
    input    			wire                             		i_cfg_acl_item_dmac_code_3_valid      , // д����Ч�ź�
					
    input    			wire [15:0]                      		i_cfg_acl_item_dmac_code_4            , // �˿�ACL����-д��dmacֵ[63:48]
    input    			wire                             		i_cfg_acl_item_dmac_code_4_valid      , // д����Ч�ź�
					
    input    			wire [15:0]                      		i_cfg_acl_item_dmac_code_5            , // �˿�ACL����-д��dmacֵ[79:64]
    input    			wire                             		i_cfg_acl_item_dmac_code_5_valid      , // д����Ч�ź�
					
    input    			wire [15:0]                      		i_cfg_acl_item_dmac_code_6            , // �˿�ACL����-д��dmacֵ[95:80]
    input    			wire                             		i_cfg_acl_item_dmac_code_6_valid      , // д����Ч�ź�
		
    // SMAC����ֵ���ã�6��16λ�ֶΣ�		
    input    			wire [15:0]                      		i_cfg_acl_item_smac_code_1            , // �˿�ACL����-д��smacֵ[15:0]
    input    			wire                             		i_cfg_acl_item_smac_code_1_valid      , // д����Ч�ź�
					
    input    			wire [15:0]                      		i_cfg_acl_item_smac_code_2            , // �˿�ACL����-д��smacֵ[31:16]
    input    			wire                             		i_cfg_acl_item_smac_code_2_valid      , // д����Ч�ź�
					
    input    			wire [15:0]                      		i_cfg_acl_item_smac_code_3            , // �˿�ACL����-д��smacֵ[47:32]
    input    			wire                             		i_cfg_acl_item_smac_code_3_valid      , // д����Ч�ź�
					
    input    			wire [15:0]                      		i_cfg_acl_item_smac_code_4            , // �˿�ACL����-д��smacֵ[63:48]
    input    			wire                             		i_cfg_acl_item_smac_code_4_valid      , // д����Ч�ź�
					
    input    			wire [15:0]                      		i_cfg_acl_item_smac_code_5            , // �˿�ACL����-д��smacֵ[79:64]
    input    			wire                             		i_cfg_acl_item_smac_code_5_valid      , // д����Ч�ź�
					
    input    			wire [15:0]                      		i_cfg_acl_item_smac_code_6            , // �˿�ACL����-д��smacֵ[95:80]
    input    			wire                             		i_cfg_acl_item_smac_code_6_valid      , // д����Ч�ź�
		
    // VLAN����ֵ���ã�4��16λ�ֶΣ�		
    input    			wire [15:0]                      		i_cfg_acl_item_vlan_code_1            , // �˿�ACL����-д��vlanֵ[15:0]
    input    			wire                             		i_cfg_acl_item_vlan_code_1_valid      , // д����Ч�ź�
					
    input    			wire [15:0]                      		i_cfg_acl_item_vlan_code_2            , // �˿�ACL����-д��vlanֵ[31:16]
    input    			wire                             		i_cfg_acl_item_vlan_code_2_valid      , // д����Ч�ź�
					
    input    			wire [15:0]                      		i_cfg_acl_item_vlan_code_3            , // �˿�ACL����-д��vlanֵ[47:32]
    input    			wire                             		i_cfg_acl_item_vlan_code_3_valid      , // д����Ч�ź�
					
    input    			wire [15:0]                      		i_cfg_acl_item_vlan_code_4            , // �˿�ACL����-д��vlanֵ[63:48]
    input    			wire                             		i_cfg_acl_item_vlan_code_4_valid      , // д����Ч�ź�

    // Ethertype����ֵ���ã�2��16λ�ֶΣ�
    input    			wire [15:0]                      		i_cfg_acl_item_ethertype_code_1       , // �˿�ACL����-д��ethertypeֵ[15:0]
    input    			wire                             		i_cfg_acl_item_ethertype_code_1_valid , // д����Ч�ź�
					
    input    			wire [15:0]                      		i_cfg_acl_item_ethertype_code_2       , // �˿�ACL����-д��ethertypeֵ[31:16]
    input    			wire                             		i_cfg_acl_item_ethertype_code_2_valid , // д����Ч�ź�

    // ACL��������
    input    			wire [7:0]                       	    i_cfg_acl_item_action_pass_state      , // �˿�ACL����-����״̬
    input    			wire                             	    i_cfg_acl_item_action_pass_state_valid, // д����Ч�ź�
				    
    input    			wire [15:0]                      	    i_cfg_acl_item_action_cb_streamhandle , // �˿�ACL����-stream_handleֵ
    input    			wire                             	    i_cfg_acl_item_action_cb_streamhandle_valid, // д����Ч�ź�
				    
    input    			wire [5:0]                       	    i_cfg_acl_item_action_flowctrl        , // �˿�ACL����-��������ѡ��
    input    			wire                             	    i_cfg_acl_item_action_flowctrl_valid  , // д����Ч�ź�
				    
    input    			wire [15:0]                      	    i_cfg_acl_item_action_txport          , // �˿�ACL����-���ķ��Ͷ˿�ӳ��
    input    			wire                             	    i_cfg_acl_item_action_txport_valid    ,  // д����Ч�ź�

    // ״̬�Ĵ���
    output             wire   [15:0]                            o_port_diag_state                  , // �˿�״̬�Ĵ�����������Ĵ�����˵������ 
    output             wire                                     o_tcam_config_busy                 , // TCAM ����æ
    output             wire                                     o_tcam_fsm_state                   , // TCAM ��ǰ״̬
    // ��ϼĴ���
    output             wire                                     o_port_rx_ultrashort_frm           , // �˿ڽ��ճ���֡(С��64�ֽ�)
    output             wire                                     o_port_rx_overlength_frm           , // �˿ڽ��ճ���֡(����MTU�ֽ�)
    output             wire                                     o_port_rx_crcerr_frm               , // �˿ڽ���CRC����֡
    output             wire  [15:0]                             o_port_rx_loopback_frm_cnt         , // �˿ڽ��ջ���֡������ֵ
    output             wire  [15:0]                             o_port_broadflow_drop_cnt          , // �˿ڽ��յ��㲥������������֡������ֵ
    output             wire  [15:0]                             o_port_multiflow_drop_cnt          , // �˿ڽ��յ��鲥������������֡������ֵ
    // ����ͳ�ƼĴ���
    output             wire  [15:0]                             o_port_rx_byte_cnt                 , // �˿�0�����ֽڸ���������ֵ
    output             wire  [15:0]                             o_port_rx_frame_cnt                  // �˿�0����֡����������ֵ  
);

/*----------- locaparameter -------*/

wire    [PORT_NUM-1:0]                  w_swlist_tx_port                    ; // ���Ͷ˿���Ϣ
wire                                    w_swlist_vld                        ; // ��Чʹ���ź�  

// rx_data_stream_cross ������������
wire                                    w_mac_port_link                     ;   
wire   [1:0]                            w_mac_port_speed                    ;         
wire                                    w_mac_port_filter_preamble_v        ;   
wire   [PORT_MNG_DATA_WIDTH-1:0]        w_mac_axi_data                      ;       
wire   [(PORT_MNG_DATA_WIDTH/8)-1:0]    w_mac_axi_data_keep                 ;        
wire                                    w_mac_axi_data_valid                ;        
wire                                    w_mac_axi_data_ready                ;             
wire                                    w_mac_axi_data_last                 ; 

// qbu �������֮���������
wire                                    w_qbu_mac_port_link                 ;   
wire   [1:0]                            w_qbu_mac_port_speed                ;         
wire                                    w_qbu_mac_port_filter_preamble_v    ;   
wire   [PORT_MNG_DATA_WIDTH-1:0]        w_qbu_mac_axi_data                  ;       
wire   [(PORT_MNG_DATA_WIDTH/8)-1:0]    w_qbu_mac_axi_data_keep             ;  
wire   [15:0]                           w_qbu_mac_axi_data_user             ;      
wire                                    w_qbu_mac_axi_data_valid            ;        
wire                                    w_qbu_mac_axi_data_ready            ;             
wire                                    w_qbu_mac_axi_data_last             ; 

// �����������������

wire                                    w_mac_time_irq                      ; // ��ʱ����ж��ź�
wire  [7:0]                             w_mac_frame_seq                     ; // ֡���к�
wire  [6:0]                             w_timestamp_addr                    ; // ��ʱ����洢�� RAM ��ַ

wire  [15:0]                            w_port_rx_byte_cnt                  ; // �˿�0�����ֽڸ���������ֵ
wire  [15:0]                            w_port_rx_frame_cnt                 ; // �˿�0����֡����������ֵ 

// wire                                    w_mac_cross_port_link               ;
wire   [1:0]                            w_mac_cross_port_speed              ;
wire   [CROSS_DATA_WIDTH-1:0]           w_mac_cross_axi_data                ;
wire   [15:0]                           w_mac_cross_axi_data_user           ;
wire   [(CROSS_DATA_WIDTH/8)-1:0]       w_mac_cross_axi_data_keep           ;
wire                                    w_mac_cross_axi_data_valid          ;
wire                                    w_mac_cross_axi_data_ready          ;
wire                                    w_mac_cross_axi_data_last           ;

wire   [CROSS_DATA_WIDTH-1:0]           w_mac_cross_port_axi_data           ; // �ӵ��ⲿ�ź�
wire   [(CROSS_DATA_WIDTH/8)-1:0]       w_mac_cross_port_axi_keep           ; // �ӵ��ⲿ�ź�
wire   [15:0]                           w_mac_cross_port_axi_user           ; // �ӵ��ⲿ�ź�
wire                                    w_mac_cross_port_axi_valid          ; // �ӵ��ⲿ�ź�
wire                                    w_mac_cross_port_axi_ready          ; // �ӵ��ⲿ�ź�
wire                                    w_mac_cross_port_axi_last           ; // �ӵ��ⲿ�ź�

// rx_frm_info_mng �������Ϣ
wire                                    w_mac_frm_info_cross_axi_data_ready ;
wire   [1:0]                            w_port_speed                        ;
wire   [2:0]                            w_vlan_pri                          ;
wire                                    w_frm_vlan_flag                     ;
wire   [PORT_NUM-1:0]                   w_rx_port                           ;
wire   [1:0]                            w_frm_cb_op                         ;
wire                                    w_frm_qbu                           ;
wire   [47:0]                           w_dmac_data                         ;
wire                                    w_damac_data_vld                    ;
wire                                    w_dmac_soc                          ;
wire                                    w_dmac_eoc                          ;
wire   [47:0]                           w_smac_data                         ;
wire                                    w_samac_data_vld                    ;
wire                                    w_smac_soc                          ;
wire                                    w_smac_eoc                          ;
wire                                    w_info_valid                        ;
wire   [11:0]                           w_vlan_id                           ;    
wire   [15:0]                           w_rtag_sequence                     ;
wire   [15:0]                           w_ethertyper                        ;

// rx_data_width output
wire   [LOOK_UP_DATA_WIDTH-1:0]         w_mac_width_port_axi_data           ;
wire                                    w_mac_width_axi_data_valid          ;

// rx_frm_acl_mng �������Ϣ
wire                                    w_mac_frm_acl_axi_data_ready        ;
wire                                    w_acl_vld                           ; 
wire    [2:0]                           w_acl_action                        ;
wire                                    w_acl_cb_frm                        ;
wire    [7:0]                           w_acl_cb_streamhandle               ;
wire    [2:0]                           w_acl_flow_ctrl                     ;
wire    [7:0]                           w_acl_forwardport                   ;
// wire                                    w_acl_find_match                    ; 
// wire   [7:0]                            w_acl_frmtype                       ; 
// wire   [15:0]                           w_acl_fetch_info                    ;
wire                                    w_acl_list_rdy_regs                 ;
 

wire   [11:0]                           w_vlanid                           ;
wire   [HASH_DATA_WIDTH - 1 : 0]        w_dmac_hash_key                    ; // Ŀ�� mac �Ĺ�ϣֵ
wire   [47 : 0]                         w_dmac                             ; // Ŀ�� mac ��ֵ
wire                                    w_dmac_hash_vld                    ; // dmac_vld
wire   [HASH_DATA_WIDTH - 1 : 0]        w_smac_hash_key                    ; // Դ mac ��ֵ��Ч��ʶ
wire   [47 : 0]                         w_smac                             ; // Դ mac ��ֵ
wire                                    w_smac_hash_vld                    ; // smac_vld

wire   [METADATA_WIDTH-1:0]             w_cross_metadata                   ; // �ۺ����� metadata ����
wire                                    w_cross_metadata_valid             ; // �ۺ����� metadata ������Ч
wire                                    w_cross_metadata_last              ; // ��Ϣ��������ʶ
wire                                    w_cross_metadata_ready             ; // ����ģ�鷴ѹ��ˮ�� 

wire   [METADATA_WIDTH-1:0]             w_cross_port_metadata              ;
wire                                    w_cross_port_metadata_valid        ;
wire                                    w_cross_port_metadata_last         ;
wire                                    w_cross_port_metadata_ready        ;

// rx_forward_mng ���ź�
wire                                    w_port_rx_ultrashort_frm           ; // �˿ڽ��ճ���֡(С��64�ֽ�)
wire                                    w_port_rx_overlength_frm           ; // �˿ڽ��ճ���֡(����MTU�ֽ�)
wire                                    w_port_rx_crcerr_frm               ; // �˿ڽ���CRC����֡
wire  [15:0]                            w_port_rx_loopback_frm_cnt         ; // �˿ڽ��ջ���֡������ֵ
wire  [15:0]                            w_port_broadflow_drop_cnt          ; // �˿ڽ��յ��㲥������������֡������ֵ
wire  [15:0]                            w_port_multiflow_drop_cnt          ; // �˿ڽ��յ��鲥������������֡������ֵ
wire  [15:0]                            w_port_diag_state                  ;  // �˿�״̬�Ĵ�����������Ĵ�����˵������ 

wire                                    w_port_rxmac_down_regs             ; // �˿ڽ��շ���MAC�ر�ʹ��
wire                                    w_port_broadcast_drop_regs         ; // �˿ڹ㲥֡����ʹ��
wire                                    w_port_multicast_drop_regs         ; // �˿��鲥֡����ʹ��
wire                                    w_port_loopback_drop_regs          ; // �˿ڻ���֡����ʹ��
wire   [47:0]                           w_port_mac_regs                    ; // �˿ڵ� MAC ��ַ
wire                                    w_port_mac_vld_regs                ; // ʹ�ܶ˿� MAC ��ַ��Ч
wire   [7:0]                            w_port_mtu_regs                    ; // MTU����ֵ
wire   [PORT_NUM-1:0]                   w_port_mirror_frwd_regs            ; // ����ת���Ĵ���������Ӧ�Ķ˿���1���򱾶˿ڽ��յ����κ�ת������֡������ת��ֵ����1�Ķ˿�
wire   [15:0]                           w_port_flowctrl_cfg_regs           ; // ������������                                                                        
wire   [4:0]                            w_port_rx_ultrashortinterval_num   ; // ֡���    

//qbu�ļĴ����ź�
wire                                    w_rx_busy                          ;
wire   [15:0]                           w_rx_fragment_cnt                  ;
wire                                    w_rx_fragment_mismatch             ;
wire   [15:0]                           w_err_rx_crc_cnt                   ;
wire   [15:0]                           w_err_rx_frame_cnt                 ;
wire   [15:0]                           w_err_fragment_cnt                 ;
wire   [15:0]                           w_rx_frames_cnt                    ;
wire   [7:0]                            w_frag_next_rx                     ; 
wire   [7:0]                            w_frame_seq                        ;

wire                                    w_verify_enabled                   ;
wire                                    w_start_verify                     ;
wire                                    w_clear_verify                     ;
wire                                    w_verify_succ                      ;
wire                                    w_verify_succ_val                  ;
wire   [7:0]                            w_verify_timer                     ;
wire                                    w_verify_timer_vld                 ;
wire   [15:0]                           w_err_verify_cnt                   ;
wire                                    w_preempt_enable                   ;

wire                                    w_dmac_vld                         ;
wire                                    w_smac_vld                         ;
wire                                    w_rtag_flag                        ; 


wire    [PORT_NUM-1:0]					w_acl_port_sel					   ;
wire									w_acl_port_sel_valid			   ;
wire									w_acl_clr_list_regs				   ;
wire	[4:0]							w_acl_item_sel_regs				   ;	

/* ------------------------------ �ڲ����������� ------------------------------- */
// assign              o_mac_cross_port_link               =      w_mac_cross_port_link        ;
assign              o_mac_cross_port_speed              =      w_mac_cross_port_speed       ;
assign              o_mac_cross_port_axi_data           =      w_mac_cross_port_axi_data    ;
assign              o_mac_cross_port_axi_user           =      w_mac_cross_port_axi_user    ;
assign              o_mac_cross_axi_data_keep           =      w_mac_cross_port_axi_keep    ;
assign              o_mac_cross_axi_data_valid          =      w_mac_cross_port_axi_valid   ;
assign              w_mac_cross_port_axi_ready          =      i_mac_cross_axi_data_ready   ;
assign              o_mac_cross_axi_data_last           =      w_mac_cross_port_axi_last    ;
  

/* ------------------------------ ����ģ������������ ------------------------------- */
// input
// assign              w_mac_port_link                     =      i_mac_port_link              ;
assign              w_mac_port_speed                    =      i_mac_port_speed             ;
assign              w_mac_port_filter_preamble_v        =      i_mac_port_filter_preamble_v ;
assign              w_mac_axi_data                      =      i_mac_axi_data               ;
assign              w_mac_axi_data_keep                 =      i_mac_axi_data_keep          ;
assign              w_mac_axi_data_valid                =      i_mac_axi_data_valid         ;
assign              o_mac_axi_data_ready                =      w_mac_axi_data_ready         ;
assign              w_mac_axi_data_last                 =      i_mac_axi_data_last          ;

assign              w_acl_port_sel                      =      i_acl_port_sel               ; 
assign 				w_acl_port_sel_valid				=	   i_acl_port_sel_valid			;  
assign              w_acl_clr_list_regs                 =      i_acl_clr_list_regs          ;   
assign              o_acl_list_rdy_regs                 =      w_acl_list_rdy_regs          ;   
assign              w_acl_item_sel_regs                 =      i_acl_item_sel_regs          ;   

assign              w_swlist_tx_port                    =      i_swlist_tx_port             ;
assign              w_swlist_vld                        =      i_swlist_vld                 ;

assign              w_port_rxmac_down_regs              =      i_port_rxmac_down_regs       ;   
assign              w_port_broadcast_drop_regs          =      i_port_broadcast_drop_regs   ;   
assign              w_port_multicast_drop_regs          =      i_port_multicast_drop_regs   ;   
assign              w_port_loopback_drop_regs           =      i_port_loopback_drop_regs    ;   
assign              w_port_mac_regs                     =      i_port_mac_regs              ;   
assign              w_port_mac_vld_regs                 =      i_port_mac_vld_regs          ;   
assign              w_port_mtu_regs                     =      i_port_mtu_regs              ;   
assign              w_port_mirror_frwd_regs             =      i_port_mirror_frwd_regs      ;   
assign              w_port_flowctrl_cfg_regs            =      i_port_flowctrl_cfg_regs     ;   
assign              w_port_rx_ultrashortinterval_num    =      i_port_rx_ultrashortinterval_num;

// output
assign              o_mac_time_irq                      =      w_mac_time_irq               ;
assign              o_mac_frame_seq                     =      w_mac_frame_seq              ;
assign              o_timestamp_addr                    =      w_timestamp_addr             ;

assign              o_port_rx_byte_cnt                  =      w_port_rx_byte_cnt           ;
assign              o_port_rx_frame_cnt                 =      w_port_rx_frame_cnt          ;

assign              o_vlan_id                           =      w_vlanid                     ;
assign              o_dmac_hash_key                     =      w_dmac_hash_key              ;
assign              o_dmac                              =      w_dmac                       ;
assign              o_dmac_vld                          =      w_dmac_vld                   ;
assign              o_smac_hash_key                     =      w_smac_hash_key              ;
assign              o_smac                              =      w_smac                       ;
assign              o_smac_vld                          =      w_smac_vld                   ;

// assign              o_rtag_flag                         =      w_rtag_flag                  ;
// assign              o_rtag_squence                      =      w_rtag_sequence              ;
// assign              o_stream_handle                     =      w_acl_cb_streamhandle        ;

assign              o_cross_metadata                    =      w_cross_port_metadata        ;
assign              o_cross_metadata_valid              =      w_cross_port_metadata_valid  ;
assign              o_cross_metadata_last               =      w_cross_port_metadata_last   ;
assign              w_cross_port_metadata_ready         =      i_cross_metadata_ready       ;

assign              o_port_rx_ultrashort_frm            =      w_port_rx_ultrashort_frm     ;
assign              o_port_rx_overlength_frm            =      w_port_rx_overlength_frm     ;   
assign              o_port_rx_crcerr_frm                =      w_port_rx_crcerr_frm         ;       
assign              o_port_rx_loopback_frm_cnt          =      w_port_rx_loopback_frm_cnt   ;   
assign              o_port_broadflow_drop_cnt           =      w_port_broadflow_drop_cnt    ;   
assign              o_port_multiflow_drop_cnt           =      w_port_multiflow_drop_cnt    ;   
assign              o_port_diag_state                   =      w_port_diag_state            ;

/* ------------------------------ ֡��ռ����ͨ· ------------------------------- */

qbu_rec #(
    .DWIDTH                           (PORT_MNG_DATA_WIDTH          ),
	.PORT_INDEX 					  (PORT_INDEX  		            )
) qbu_rec_inst (          
    .i_clk                            (i_clk                        ),
    .i_rst                            (i_rst                        ),
    //�ӿڲ�����������
    .i_mac_port_speed                 (w_mac_port_speed             ),
    .i_mac_axi_data                   (w_mac_axi_data               ), 
    .i_mac_axi_data_keep              (w_mac_axi_data_keep          ), 
    .i_mac_axi_data_valid             (w_mac_axi_data_valid         ), 
    .o_mac_axi_data_ready             (w_mac_axi_data_ready         ), 
    .i_mac_axi_data_last              (w_mac_axi_data_last          ), 
    //�����tx_mac����֤qbu����
    .o_qbu_verify_valid               (i_qbu_verify_valid           ),
    .o_qbu_response_valid             (i_qbu_response_valid         ),
    //���qbu emac��pmacͨ�����ݣ�emacͨ�������ж����
    .o_qbu_rx_axis_portspeed          (w_qbu_mac_port_speed         ),
    .o_qbu_rx_axis_data               (w_qbu_mac_axi_data           ),
    .o_qbu_rx_axis_user               (w_qbu_mac_axi_data_user      ),
    .o_qbu_rx_axis_keep               (w_qbu_mac_axi_data_keep      ),
    .o_qbu_rx_axis_last               (w_qbu_mac_axi_data_last      ),
    .o_qbu_rx_axis_valid              (w_qbu_mac_axi_data_valid     ),
    .i_qbu_rx_axis_ready              (w_qbu_mac_axi_data_ready     ),  

    .o_dmac			                  (w_dmac_data                  ),      
    .o_smac 			              (w_smac_data                  ),          
    // .o_port_speed                     (w_port_speed                 ),      
    .o_vlan_pri                       (w_vlan_pri                   ),      
    .o_vlan_id                        (w_vlan_id                    ),      
    .o_frm_vlan_flag                  (w_frm_vlan_flag              ),      
    .o_frm_qbu                        (w_frm_qbu                    ),      
    .o_frm_discard                    (w_frm_discard                ),      
    .o_rtag_sequence                  (w_rtag_sequence              ),      
    .o_rtag_flag                      (w_rtag_flag                  ),      
    .o_ethertype 	                  (w_ethertyper                 ),      
    .o_info_valid                     (w_info_valid                 ),      
    // // ��ʱ����ź�
    .o_mac_time_irq                   (w_mac_time_irq               ),  
    .o_mac_frame_seq                  (w_mac_frame_seq              ),  
    .o_timestamp_addr                 (w_timestamp_addr             ),     
    //qbu�Ĵ�������
    .i_default_vlan_id                (12'd0 ), // �ȴ�����߼�
    .i_default_vlan_pri               (3'd0  ), // �ȴ�����߼�
    .i_default_vlan_valid             (1'd0  ), // �ȴ�����߼�

    .i_verify_enabled	              (w_verify_enabled	            ),
    .i_verify_timer		              (w_verify_timer		        ),
    .i_verify_timer_valid             (w_verify_timer_valid         ),
    .i_reset 			              (w_reset 			            ),
    .i_start_verify     	          (w_start_verify               ),
    .i_clear_verify     	          (w_clear_verify               ),
    
    .o_rx_busy                        (w_rx_busy             	    ), 
    .o_rx_fragment_cnt                (w_rx_fragment_cnt     	    ), 
    .o_rx_fragment_mismatch           (w_rx_fragment_mismatch	    ), 
    .o_err_rx_crc_cnt                 (w_err_rx_crc_cnt      	    ), 
    .o_err_rx_frame_cnt               (w_err_rx_frame_cnt    	    ), 
    .o_err_fragment_cnt               (w_err_fragment_cnt    	    ), 
    .o_rx_frames_cnt                  (w_rx_frames_cnt       	    ), 
    .o_frag_next_rx                   (w_frag_next_rx        	    ), 
    .o_err_verify_cnt                 (w_err_verify_cnt             ),
    .o_preempt_enable                 (w_preempt_enable             ),
    .o_frame_seq                      (w_frame_seq           	    )  
);

/* ----------------------------- ������������Ϣ��ȡ����ˮ�߲����� -------------------------------- */

// rx_frm_info_mng#(
//     .PORT_NUM                       ( PORT_NUM                       )   ,
//     .PORT_MNG_DATA_WIDTH            ( PORT_MNG_DATA_WIDTH            )   ,
//     .CROSS_DATA_WIDTH               ( CROSS_DATA_WIDTH               )   ,
//     .PORT_INDEX                     ( PORT_INDEX                     )
// )rx_frm_info_mng_inst (
//     .i_clk                          ( i_clk                          )   ,
//     .i_rst                          ( i_rst                          )   ,
//     /*---------------------------------------- �� PORT �ۺ������� ----------------------------------*/
//     // .i_mac_port_link                ( w_qbu_mac_port_link            )   ,
//     .i_mac_port_speed               ( w_qbu_mac_port_speed           )   ,
//     .i_mac_port_axi_data            ( w_qbu_mac_axi_data             )   ,
//     .i_mac_axi_data_keep            ( w_qbu_mac_axi_data_keep        )   ,
//     .i_mac_axi_data_user            ( w_qbu_mac_axi_data_user        )   ,  
//     .i_mac_axi_data_valid           ( w_qbu_mac_axi_data_valid       )   ,
//     .o_mac_axi_data_ready           ( w_qbu_mac_axi_data_ready       )   ,
//     .i_mac_axi_data_last            ( w_qbu_mac_axi_data_last        )   ,
//     // �Ĵ�����������
//     .i_default_vlan_id              (12'd0 ), // �ȴ�����߼�
//     .i_default_vlan_pri             (3'd0  ), // �ȴ�����߼�
//     .i_default_vlan_valid           (1'd0  ), // �ȴ�����߼�

//     /* �� PORT ������Ϣ�� */
//     .o_port_speed                   ( w_port_speed                   )   ,
//     .o_vlan_pri                     ( w_vlan_pri                     )   ,
//     .o_frm_vlan_flag                ( w_frm_vlan_flag                )   ,
//     .o_rx_port                      ( w_rx_port                      )   ,
//     .o_frm_qbu                      ( w_frm_qbu                      )   ,
//     .o_frm_discard                  ( w_frm_discard                  )   ,  
//     .o_vlan_id                      ( w_vlan_id                      )   ,  
//     .o_rtag_sequence                ( w_rtag_sequence                )   ,  
//     .o_ethertyper                   ( w_ethertyper                   )   ,  
//     /*-------------------------- �ڲ������������Ϣ�� ----------------------------*/
//     .o_dmac_data                    ( w_dmac_data                    )   ,
//     .o_damac_data_vld               ( w_damac_data_vld               )   ,
//     .o_dmac_soc                     ( w_dmac_soc                     )   ,
//     .o_dmac_eoc                     ( w_dmac_eoc                     )   ,
//     .o_smac_data                    ( w_smac_data                    )   ,
//     .o_samac_data_vld               ( w_samac_data_vld               )   ,
//     .o_smac_soc                     ( w_smac_soc                     )   ,
//     .o_smac_eoc                     ( w_smac_eoc                     )   ,
//     .o_frm_info_vld                 ( w_frm_info_vld                 )   ,
//     .o_broadcast_frm_en             ( w_broadcast_frm_en             )   ,
//     .o_multicast_frm_en             ( w_multicast_frm_en             )   ,
//     .o_flood_frm_en                 ( w_flood_frm_en                 )
// );

// --------------- �����Ҫ������ 144bit
// rx_data_width #(
//     .INPUT_WIDTH                    ( PORT_MNG_DATA_WIDTH           ),
//     .OUTPUT_WIDTH                   ( LOOK_UP_DATA_WIDTH            )
// ) rx_data_width_inst (
//     .i_clk                          ( i_clk                         ),
//     .i_rst                          ( i_rst                         ),
//     .i_mac_port_filter_preamble_v   ( i_mac_port_filter_preamble_v  ),
//     .i_mac_axi_data                 ( w_qbu_mac_axi_data            ),
//     .i_mac_axi_data_keep            ( w_qbu_mac_axi_data_keep       ),
//     .i_mac_axi_data_valid           ( w_qbu_mac_axi_data_valid      ),
//     .o_mac_axi_data_ready           (                               ),
//     .i_mac_axi_data_last            ( w_qbu_mac_axi_data_last       ),

//     .o_mac_cross_port_axi_data      ( w_mac_width_port_axi_data     ),
//     .o_mac_cross_axi_data_valid     ( w_mac_width_axi_data_valid    )
// );

rx_acllookup_data rx_acllookup_data_inst (
    .i_clk                          ( i_clk                         ),
    .i_rst                          ( i_rst                         ),

    .i_dmac_data                    ( w_dmac_data                   ), 
    .i_smac_data                    ( w_smac_data                   ), 

    .i_vlan_id                      ( w_vlan_id                     ),
    .i_vlan_pri                     ( w_vlan_pri                    ),
    .i_ethertyper                   ( w_ethertyper                  ),
    .i_info_vld                     ( w_info_valid                  ),

    .o_mac_cross_port_axi_data      ( w_mac_width_port_axi_data     ),
    .o_mac_cross_axi_data_valid     ( w_mac_width_axi_data_valid    )
);

// --------------

//tcam_top #(
//    .LOOK_UP_DATA_WIDTH             ( LOOK_UP_DATA_WIDTH          ),   // ��Ҫ��ѯ��������λ��
//    .REG_ADDR_BUS_WIDTH             ( REG_ADDR_BUS_WIDTH          ),   // ���� MAC ������üĴ�����ַλ��
//    .REG_DATA_BUS_WIDTH             ( REG_DATA_BUS_WIDTH          ),   // ���� MAC ������üĴ�������λ��
//    .ACTION_WIDTH                   ( 24                          ),   // ACTION
//    .CAM_NUM                        ( 256                         )    // ��������
//) tcam_top_inst (           
//    .i_clk                          ( i_clk                       ),
//    .i_rst                          ( i_rst                       ),
//    /*---------------------------------------- ƥ���������� ------------------------------------------*/
//    .i_look_up_data                 ( w_mac_width_port_axi_data   ),
//    .i_look_up_data_vld             ( w_mac_width_axi_data_valid  ),
//    /*---------------------------------------- ƥ�� ACTION ��� --------------------------------------*/
//    // .o_acl_frmtype                  ( w_acl_frmtype               ),
//    // .o_acl_fetchinfo                ( w_acl_fetch_info            ),
//    .o_acl_action                   ( w_acl_action                ),
//    .o_acl_cb_frm                   ( w_acl_cb_frm                ),
//    .o_acl_cb_streamhandle          ( w_acl_cb_streamhandle       ),
//    .o_acl_flow_ctrl                ( w_acl_flow_ctrl             ),
//    .o_acl_forwardport              ( w_acl_forwardport           ),  
//    .o_acl_vld                      ( w_acl_vld                   ),
//    /*---------------------------------------- �Ĵ������ýӿ� -----------------------------------------*/
//    .o_tcam_busy                    ( o_tcam_config_busy          ) // ������ϲ��������tcam��busy
//    // �Ĵ��������ź�       
//    //.i_refresh_list_pulse           ( i_refresh_list_pulse        ), // ˢ�¼Ĵ����б�״̬�Ĵ����Ϳ��ƼĴ�����
//    //.i_switch_err_cnt_clr           ( i_switch_err_cnt_clr        ), // ˢ�´��������
//    //.i_switch_err_cnt_stat          ( i_switch_err_cnt_stat       ), // ˢ�´���״̬�Ĵ���
//    // �Ĵ���д���ƽӿ�       
//    //.i_switch_reg_bus_we            ( i_switch_reg_bus_we         ), // �Ĵ���дʹ��
//    //.i_switch_reg_bus_we_addr       ( i_switch_reg_bus_we_addr    ), // �Ĵ���д��ַ
//    //.i_switch_reg_bus_we_din        ( i_switch_reg_bus_we_din     ), // �Ĵ���д����
//    //.i_switch_reg_bus_we_din_v      ( i_switch_reg_bus_we_din_v   ), // �Ĵ���д����ʹ��
//    // �Ĵ��������ƽӿ�       
//    //.i_switch_reg_bus_rd            ( i_switch_reg_bus_rd         ), // �Ĵ�����ʹ��
//    //.i_switch_reg_bus_rd_addr       ( i_switch_reg_bus_rd_addr    ), // �Ĵ�������ַ
//    //.o_switch_reg_bus_we_dout       ( o_switch_reg_bus_we_dout    ), // �����Ĵ�������
//    //.o_switch_reg_bus_we_dout_v     ( o_switch_reg_bus_we_dout_v  )  // ��������Чʹ��
//  );


tcam_top #(
	 .LOOK_UP_DATA_WIDTH             ( LOOK_UP_DATA_WIDTH    ),
	 .PORT_MNG_DATA_WIDTH            ( PORT_MNG_DATA_WIDTH   ),
	 .REG_ADDR_BUS_WIDTH             ( REG_ADDR_BUS_WIDTH    ),
	 .REG_DATA_BUS_WIDTH             ( REG_DATA_BUS_WIDTH    ),
	 .PORT_ID                        ( PORT_INDEX            ),
	 .CAM_NUM                        ( CAM_NUM               )
) tcam_top_inst (
	 .i_clk                          ( i_clk                        	 ),
	 .i_rst                          ( i_rst                        	 ),
	 //
	 .i_look_up_data                 ( w_mac_width_port_axi_data     	 ),
	 .i_look_up_data_vld             ( w_mac_width_axi_data_valid    	 ),
	 
	 .o_acl_action                   ( w_acl_action               		 ),
	 .o_acl_cb_frm                   ( w_acl_cb_frm               		 ),
	 .o_acl_cb_streamhandle          ( w_acl_cb_streamhandle      		 ),
	 .o_acl_flow_ctrl                ( w_acl_flow_ctrl            		 ),
	 .o_acl_forwardport              ( w_acl_forwardport          		 ),
	 .o_acl_vld                      ( w_acl_vld                  		 ),
	 .o_tcam_busy                    ( o_tcam_config_busy                ),
	 
	 // New configuration interface
	 .i_cfg_acl_port_sel             ( w_acl_port_sel       		),   //
	 .i_cfg_acl_port_sel_valid       ( w_acl_port_sel_valid       	),   //
	 .i_cfg_acl_clr_list_regs        ( w_acl_clr_list_regs        	),   //
	 .o_cfg_acl_list_rdy_regs        ( w_acl_list_rdy_regs        	),   //
	 .o_cfg_acl_clr_busy_regs		 (),

	 // DMAC
	 .i_cfg_acl_item_dmac_code_1     	(i_cfg_acl_item_dmac_code_1     ),  
	 .i_cfg_acl_item_dmac_code_1_valid	(i_cfg_acl_item_dmac_code_1_valid),
	 .i_cfg_acl_item_dmac_code_2     	(i_cfg_acl_item_dmac_code_2     ),  
	 .i_cfg_acl_item_dmac_code_2_valid	(i_cfg_acl_item_dmac_code_2_valid),
	 .i_cfg_acl_item_dmac_code_3     	(i_cfg_acl_item_dmac_code_3     ),  
	 .i_cfg_acl_item_dmac_code_3_valid	(i_cfg_acl_item_dmac_code_3_valid),
	 .i_cfg_acl_item_dmac_code_4     	(i_cfg_acl_item_dmac_code_4     ),  
	 .i_cfg_acl_item_dmac_code_4_valid	(i_cfg_acl_item_dmac_code_4_valid),
	 .i_cfg_acl_item_dmac_code_5     	(i_cfg_acl_item_dmac_code_5     ),  
	 .i_cfg_acl_item_dmac_code_5_valid	(i_cfg_acl_item_dmac_code_5_valid),
	 .i_cfg_acl_item_dmac_code_6     	(i_cfg_acl_item_dmac_code_6     ),  
	 .i_cfg_acl_item_dmac_code_6_valid	(i_cfg_acl_item_dmac_code_6_valid),
																		
	 // SMAC                                       
	 .i_cfg_acl_item_smac_code_1     	(i_cfg_acl_item_smac_code_1     ),       
	 .i_cfg_acl_item_smac_code_1_valid	(i_cfg_acl_item_smac_code_1_valid),
	 .i_cfg_acl_item_smac_code_2     	(i_cfg_acl_item_smac_code_2     ),       
	 .i_cfg_acl_item_smac_code_2_valid	(i_cfg_acl_item_smac_code_2_valid),
	 .i_cfg_acl_item_smac_code_3     	(i_cfg_acl_item_smac_code_3     ),
	 .i_cfg_acl_item_smac_code_3_valid	(i_cfg_acl_item_smac_code_3_valid),
	 .i_cfg_acl_item_smac_code_4     	(i_cfg_acl_item_smac_code_4     ),
	 .i_cfg_acl_item_smac_code_4_valid	(i_cfg_acl_item_smac_code_4_valid),
	 .i_cfg_acl_item_smac_code_5     	(i_cfg_acl_item_smac_code_5     ),
	 .i_cfg_acl_item_smac_code_5_valid	(i_cfg_acl_item_smac_code_5_valid),
	 .i_cfg_acl_item_smac_code_6     	(i_cfg_acl_item_smac_code_6     ),
	 .i_cfg_acl_item_smac_code_6_valid	(i_cfg_acl_item_smac_code_6_valid),

	 // VLAN
	 .i_cfg_acl_item_vlan_code_1     	(i_cfg_acl_item_vlan_code_1     ),
	 .i_cfg_acl_item_vlan_code_1_valid	(i_cfg_acl_item_vlan_code_1_valid),
	 .i_cfg_acl_item_vlan_code_2     	(i_cfg_acl_item_vlan_code_2     ),
	 .i_cfg_acl_item_vlan_code_2_valid	(i_cfg_acl_item_vlan_code_2_valid),
	 .i_cfg_acl_item_vlan_code_3     	(i_cfg_acl_item_vlan_code_3     ),
	 .i_cfg_acl_item_vlan_code_3_valid	(i_cfg_acl_item_vlan_code_3_valid),
	 .i_cfg_acl_item_vlan_code_4     	(i_cfg_acl_item_vlan_code_4     ),
	 .i_cfg_acl_item_vlan_code_4_valid	(i_cfg_acl_item_vlan_code_4_valid),

	 // Ethertype
	 .i_cfg_acl_item_ethertype_code_1					(i_cfg_acl_item_ethertype_code_1		),
	 .i_cfg_acl_item_ethertype_code_1_valid				(i_cfg_acl_item_ethertype_code_1_valid	),
	 .i_cfg_acl_item_ethertype_code_2					(i_cfg_acl_item_ethertype_code_2		),
	 .i_cfg_acl_item_ethertype_code_2_valid				(i_cfg_acl_item_ethertype_code_2_valid	),
														
	 // Action                                           
	 .i_cfg_acl_item_action_pass_state					(i_cfg_acl_item_action_pass_state				),
	 .i_cfg_acl_item_action_pass_state_valid			(i_cfg_acl_item_action_pass_state_valid		),
	 .i_cfg_acl_item_action_cb_streamhandle				(i_cfg_acl_item_action_cb_streamhandle			),
	 .i_cfg_acl_item_action_cb_streamhandle_valid		(i_cfg_acl_item_action_cb_streamhandle_valid	),
	 .i_cfg_acl_item_action_flowctrl 					(i_cfg_acl_item_action_flowctrl 				),
	 .i_cfg_acl_item_action_flowctrl_valid				(i_cfg_acl_item_action_flowctrl_valid			),
	 .i_cfg_acl_item_action_txport   					(i_cfg_acl_item_action_txport   				),
	 .i_cfg_acl_item_action_txport_valid				(i_cfg_acl_item_action_txport_valid			),

	 .w_action_wea                   			    () 
	 // .o_fsm_state                    (w_fsm_state) // Removed in tcam_top? Let's check.
	 // Checking tcam_top.v again... it has w_fsm_state output?
	 // tcam_top.v: output wire [3:0] w_fsm_state
	 // Wait, I need to check if I missed it in my read.
	 // Yes, line 323: wire [3:0] w_fsm_state; but is it an output port?
	 // In tcam_top module definition:
	 // output w_action_wea,
	 // ...
	 // output wire o_tcam_busy,
	 // ...
	 // It doesn't seem to have w_fsm_state as a port in the module declaration I read earlier.
	 // Let me re-read the module declaration part of tcam_top.v carefully.
);



rx_mac_hash_calc#(
    .CWIDTH                         ( HASH_DATA_WIDTH                )
)rx_mac_hash_calc_inst (           
    .i_clk                          ( i_clk                          )    ,   // 250MHz
    .i_rst                          ( i_rst                          )    ,
    /*---------------------------------------- �Ĵ������ýӿ� -------------------------------------------*/
    .i_hash_poly_regs               ( i_hash_ploy_regs               )    ,
    .i_hash_init_val_regs           ( i_hash_init_val_regs           )    ,
    .i_hash_regs_vld                ( i_hash_regs_vld                )    ,
    /*--------------------------------- ��Ϣ��ȡģ������� MAC ��Ϣ -------------------------------------*/
    .i_vlan_id                      ( w_vlan_id                      )    ,
    .i_dmac_data                    ( w_dmac_data                    )    , // Ŀ�� MAC ��ַ��ֵ
    .i_dmac_data_vld                ( w_info_valid                   )    , // ������Чֵ 
    .i_smac_data                    ( w_smac_data                    )    , // Դ MAC ��ַ��ֵ
    .i_smac_data_vld                ( w_info_valid                   )    , // ������Чֵ 
    /*--------------------------------- ��� hash �ļ����� -------------------------------------*/     
    .o_vlan_id                      ( w_vlanid                       )    ,
    .o_dmac_hash_key                ( w_dmac_hash_key                )    ,
    .o_dmac                         ( w_dmac                         )    ,
    .o_dmac_hash_vld                ( w_dmac_vld                     )    ,
    .o_smac_hash_key                ( w_smac_hash_key                )    ,
    .o_smac                         ( w_smac                         )    ,
    .o_smac_hash_vld                ( w_smac_vld                     )            
);

rx_forward_mng#(
    .PORT_NUM                           ( PORT_NUM                       ) ,
    .PORT_MNG_DATA_WIDTH                ( PORT_MNG_DATA_WIDTH            ) ,
    .METADATA_WIDTH                     ( METADATA_WIDTH                 ) ,
    .PORT_INDEX                         ( PORT_INDEX                     ) ,
    .CROSS_DATA_WIDTH                   ( CROSS_DATA_WIDTH               )
)rx_forward_mng_inst (
    .i_clk                              ( i_clk                          ) ,
    .i_rst                              ( i_rst                          ) ,
    /* ����ת����صļĴ��� */
    .i_port_rxmac_down_regs             ( w_port_rxmac_down_regs         ) ,
    .i_port_broadcast_drop_regs         ( w_port_broadcast_drop_regs     ) ,
    .i_port_multicast_drop_regs         ( w_port_multicast_drop_regs     ) ,
    .i_port_loopback_drop_regs          ( w_port_loopback_drop_regs      ) ,
    .i_port_mac_regs                    ( w_port_mac_regs                ) ,
    .i_port_mac_vld_regs                ( w_port_mac_vld_regs            ) ,
    .i_port_mtu_regs                    ( w_port_mtu_regs                ) ,
    .i_port_mirror_frwd_regs            ( w_port_mirror_frwd_regs        ) ,
    .i_port_flowctrl_cfg_regs           (16'h00),//( w_port_flowctrl_cfg_regs       ) ,
    .i_port_rx_ultrashortinterval_num   ( w_port_rx_ultrashortinterval_num) ,
    /* rx_frm_info_mng input ����Ϣ�� */
    .i_rtag_flag                        ( w_rtag_flag                    ) ,
    .i_ethertype                        ( w_ethertyper                   ) ,
    .i_rtag_sequence                    ( w_rtag_sequence                ) ,  
    .i_port_speed                       ( w_qbu_mac_port_speed           ) ,
    .i_vlan_pri                         ( w_vlan_pri                     ) ,
    .i_frm_vlan_flag                    ( w_frm_vlan_flag                ) ,
    // .i_rx_port                          ( w_rx_port                      ) ,
    .i_frm_discard                      ( w_frm_discard                  ) ,  
    .i_frm_qbu                          ( w_frm_qbu                      ) ,
    .i_timestamp_addr                   ( w_timestamp_addr               ) ,
    .i_info_valid                       ( w_info_valid                   ) ,
    /* ���ģ����ݹ�ϣֵ���صļ����� */
    .i_swlist_port_broadcast            (i_swlist_port_broadcast         ) ,
    .i_swlist_tx_port                   ( w_swlist_tx_port               ) ,
    .i_swlist_vld                       ( w_swlist_vld                   ) ,
    /* ACL ƥ���������ֶ� */
    .i_acl_vld                          ( w_acl_vld                      ) ,
    .i_acl_action                       ( w_acl_action                   ) ,
    .i_acl_cb_frm                       ( w_acl_cb_frm                   ) ,
    .i_acl_cb_streamhandle              ( w_acl_cb_streamhandle          ) ,
    .i_acl_flow_ctrl                    ( w_acl_flow_ctrl                ) ,
    .i_acl_forwardport                  ( w_acl_forwardport              ) ,  
    // .i_acl_find_match                   ( w_acl_find_match               ) ,
    // .i_acl_frmtype                      ( w_acl_frmtype                  ) ,
    // .i_acl_fetch_info                   ( w_acl_fetch_info               ) ,
    // .i_frm_cb_op                        ( w_frm_cb_op                    ) ,
    /* �� PORT �ۺ����������� */
    .i_mac_port_axi_data                ( w_qbu_mac_axi_data             ) ,
    .i_mac_axi_data_user                ( w_qbu_mac_axi_data_user        ) ,
    .i_mac_axi_data_keep                ( w_qbu_mac_axi_data_keep        ) ,
    .i_mac_axi_data_valid               ( w_qbu_mac_axi_data_valid       ) ,
    .o_mac_axi_data_ready               ( w_qbu_mac_axi_data_ready       ) ,  
    .i_mac_axi_data_last                ( w_qbu_mac_axi_data_last        ) ,
    /* �� PORT �ۺ���������� */
    .o_mac_port_axi_data                ( w_mac_cross_axi_data           ) ,
    .o_mac_axi_data_user                ( w_mac_cross_axi_data_user      ) ,
    .o_mac_axi_data_keep                ( w_mac_cross_axi_data_keep      ) ,
    .o_mac_axi_data_valid               ( w_mac_cross_axi_data_valid     ) ,
    .i_mac_axi_data_ready               ( w_mac_cross_axi_data_ready     ) ,
    .o_mac_axi_data_last                ( w_mac_cross_axi_data_last      ) ,
    /* �� PORT �ۺ���Ϣ�� */
    .o_cross_metadata                   ( w_cross_metadata               ) ,
    .o_cross_metadata_valid             ( w_cross_metadata_valid         ) ,
    .o_cross_metadata_last              ( w_cross_metadata_last          ) ,
    .i_cross_metadata_ready             ( w_cross_metadata_ready         ) ,
    /* ��ϼĴ��� */
    .o_port_rx_ultrashort_frm           ( w_port_rx_ultrashort_frm       ) ,
    .o_port_rx_overlength_frm           ( w_port_rx_overlength_frm       ) ,
    .o_port_rx_crcerr_frm               ( w_port_rx_crcerr_frm           ) ,
    .o_port_rx_loopback_frm_cnt         ( w_port_rx_loopback_frm_cnt     ) ,
    .o_port_broadflow_drop_cnt          ( w_port_broadflow_drop_cnt      ) ,
    .o_port_multiflow_drop_cnt          ( w_port_multiflow_drop_cnt      ) ,
    .o_port_diag_state                  ( w_port_diag_state              )
);


rx_port_cache_mng#(
    .PORT_NUM                           (PORT_NUM                               ),        // �������Ķ˿���
    .PORT_MNG_DATA_WIDTH                (PORT_MNG_DATA_WIDTH                    ),        // Mac_port_mng ����λ��
    .METADATA_WIDTH                     (METADATA_WIDTH                         ),        // ��Ϣ��λ��
    .CROSS_DATA_WIDTH                   (CROSS_DATA_WIDTH                       ),        // �ۺ��������
    .PORT_FIFO_PRI_NUM                  (PORT_FIFO_PRI_NUM                      ),        // ���ȼ�FIFO����
    .RAM_DEPTH                          (1024                                   ),        // RAM���
    .RAM_ADDR_WIDTH                     (10                                     ),        // RAM��ַ���
    .FIFO_DEPTH                         (512                                    ),        // FIFO���
    .REQ_TIMEOUT_CNT                    (1250                                   ),        // req��ʱ����ֵ(5us @ 250MHz)
    .TIMEOUT_CNT_WIDTH                  (11                                     )         // ��ʱ������λ��
)rx_port_cache_mng_inst0 (
    .i_clk                              (i_clk                                  ),        // 250MHz
    .i_rst                              (i_rst                                  ),
    /*---------------------------------------- �����MAC������ -------------------------------------------*/
    .i_mac_axi_data                     ( w_mac_cross_axi_data                  ),        // �˿�������
    .i_mac_axi_data_keep                ( w_mac_cross_axi_data_keep             ),        // �˿����������룬��Ч�ֽ�ָʾ
    .i_mac_axi_data_valid               ( w_mac_cross_axi_data_valid            ),        // �˿�������Ч
    .o_mac_axi_data_ready               ( w_mac_cross_axi_data_ready            ),        // �˿����ݾ����ź�,��ʾ��ǰģ��׼���ý�������
    .i_mac_axi_data_last                ( w_mac_cross_axi_data_last             ),        // ������������ʶ
    .i_mac_axi_data_user                ( w_mac_cross_axi_data_user             ),        // ֡������Ϣ
    /*---------------------------------------- �����metadata�� -------------------------------------------*/
    .i_cross_metadata                   ( w_cross_metadata                      ),        // ����metadata����
    .i_cross_metadata_valid             ( w_cross_metadata_valid                ),        // ����metadata������Ч�ź�
    .i_cross_metadata_last              ( w_cross_metadata_last                 ),        // ����metadata������ʶ
    .o_cross_metadata_ready             ( w_cross_metadata_ready                ),        // metadata��ѹ��ˮ��
    /*---------------------------------------- ������������ߵ������� -------------------------------------------*/
    .o_mac_cross_port_axi_data          (w_mac_cross_port_axi_data              ),        // �˿������������λ��ʾcrcerr
    .o_mac_cross_port_axi_user          (w_mac_cross_port_axi_user              ),
    .o_mac_cross_axi_data_keep          (w_mac_cross_port_axi_keep              ),        // �˿����������룬��Ч�ֽ�ָʾ
    .o_mac_cross_axi_data_valid         (w_mac_cross_port_axi_valid             ),        // �˿�������Ч
    .i_mac_cross_axi_data_ready         (w_mac_cross_port_axi_ready             ),        // �������߾ۺϼܹ���ѹ��ˮ���ź�
    .o_mac_cross_axi_data_last          (w_mac_cross_port_axi_last              ),        // ������������ʶ
    /*---------------------------------------- ������������ߵ�metadata�� -------------------------------------------*/
    .o_cross_metadata                   (w_cross_port_metadata                  ),        // �ۺ�����metadata����
    .o_cross_metadata_valid             (w_cross_port_metadata_valid            ),        // �ۺ�����metadata������Ч�ź�
    .o_cross_metadata_last              (w_cross_port_metadata_last             ),        // ��Ϣ��������ʶ
    .i_cross_metadata_ready             (w_cross_port_metadata_ready            ),        // ����ģ�鷴ѹ��ˮ��
     
    /*---------------------------------------- �� PORT �ؼ�֡�ۺ���Ϣ�� -------------------------------------------*/
    .o_emac_port_axi_data               (o_emac_port_axi_data                   ) , // �˿������������λ��ʾcrcerr
    .o_emac_port_axi_user               (o_emac_port_axi_user                   ) ,
    .o_emac_axi_data_keep               (o_emac_axi_data_keep                   ) , // �˿����������룬��Ч�ֽ�ָʾ
    .o_emac_axi_data_valid              (o_emac_axi_data_valid                  ) , // �˿�������Ч
    .i_emac_axi_data_ready              (i_emac_axi_data_ready                  ) , // �������߾ۺϼܹ���ѹ��ˮ���ź�
    .o_emac_axi_data_last               (o_emac_axi_data_last                   ) , // ������������ʶ 
    .o_emac_metadata                    (o_emac_metadata                        ) , // ���� metadata ����
    .o_emac_metadata_valid              (o_emac_metadata_valid                  ) , // ���� metadata ������Ч�ź�
    .o_emac_metadata_last               (o_emac_metadata_last                   ) , // ��Ϣ��������ʶ
    .i_emac_metadata_ready              (i_emac_metadata_ready                  ) , // ����ģ�鷴ѹ��ˮ�� 
    /*---------------------------------------- �뷢�Ͷ˵�req-ack���� / CB -------------------------------------------*/
    .i_pass_en                          (i_pass_en                              ),        // �жϽ�������Խ��ո�֡
    .i_discard_en                       (i_discard_en                           ),        // �жϽ�������Զ�����֡
    .i_judge_finish                     (i_judge_finish                         ),        // �жϽ������ʾ���α��ĵ��ж����
                     
    .o_rtag_flag                        (o_rtag_flag                            ),        // ���rtag flag�����Ͷ�
    .o_rtag_squence                     (o_rtag_squence                         ),        // ���rtag flag�����Ͷ�
    .o_stream_handle                    (o_stream_handle                        ),        // ���rtag flag�����Ͷ�

    .o_tx_req                           (o_tx_req                               ),        // ���Ͷ˵�req�ź�
    .i_mac_tx0_ack                      (i_mac_tx0_ack                          ),        // �˿�0��Ӧʹ���ź�
    .i_mac_tx0_ack_rst                  (i_mac_tx0_ack_rst                      ),        // �˿�0���ȼ��������
    .i_mac_tx1_ack                      (i_mac_tx1_ack                          ),        // �˿�1��Ӧʹ���ź�
    .i_mac_tx1_ack_rst                  (i_mac_tx1_ack_rst                      ),        // �˿�1���ȼ��������
    .i_mac_tx2_ack                      (i_mac_tx2_ack                          ),        // �˿�2��Ӧʹ���ź�
    .i_mac_tx2_ack_rst                  (i_mac_tx2_ack_rst                      ),        // �˿�2���ȼ��������
    .i_mac_tx3_ack                      (i_mac_tx3_ack                          ),        // �˿�3��Ӧʹ���ź�
    .i_mac_tx3_ack_rst                  (i_mac_tx3_ack_rst                      ),        // �˿�3���ȼ��������
    .i_mac_tx4_ack                      (i_mac_tx4_ack                          ),        // �˿�4��Ӧʹ���ź�
    .i_mac_tx4_ack_rst                  (i_mac_tx4_ack_rst                      ),        // �˿�4���ȼ��������
    .i_mac_tx5_ack                      (i_mac_tx5_ack                          ),        // �˿�5��Ӧʹ���ź�
    .i_mac_tx5_ack_rst                  (i_mac_tx5_ack_rst                      ),        // �˿�5���ȼ��������
    .i_mac_tx6_ack                      (i_mac_tx6_ack                          ),        // �˿�6��Ӧʹ���ź�
    .i_mac_tx6_ack_rst                  (i_mac_tx6_ack_rst                      ),        // �˿�6���ȼ��������
    .i_mac_tx7_ack                      (i_mac_tx7_ack                          ),        // �˿�7��Ӧʹ���ź�
    .i_mac_tx7_ack_rst                  (i_mac_tx7_ack_rst                      ),        // �˿�7���ȼ��������
    /*---------------------------------------- ƽ̨�Ĵ������� -------------------------------------------*/
    .i_port_rxmac_down_regs             (1'b0                                   ),        // �˿ڽ��շ���MAC�ر�ʹ��
    .i_port_broadcast_drop_regs         (1'b0                                   ),        // �˿ڹ㲥֡����ʹ��
    .i_port_multicast_drop_regs         (1'b0                                   ),        // �˿��鲥֡����ʹ��
    .i_port_loopback_drop_regs          (1'b0                                   ),        // �˿ڻ���֡����ʹ��
    .i_port_mac_regs                    (48'h0                                  ),        // �˿ڵ�MAC��ַ
    .i_port_mac_vld_regs                (1'b0                                   ),        // ʹ�ܶ˿�MAC��ַ��Ч
    .i_port_mtu_regs                    (16'd1518                               ),        // MTU����ֵ
    .i_port_mirror_frwd_regs            ({PORT_NUM{1'b0}}                       ),        // ����ת���Ĵ���
    .i_port_flowctrl_cfg_regs           (32'h0                                  ),        // ������������
    .i_port_rx_ultrashortinterval_num   (16'd64                                 ),        // ֡���
    /*---------------------------------------- ACL�Ĵ��� -------------------------------------------*/
    .i_acl_port_sel                     (3'b0                                   ),        // ѡ��Ҫ���õĶ˿�
    .i_acl_clr_list_regs                (1'b0                                   ),        // ��ռĴ����б�
    .o_acl_list_rdy_regs                (                                       ),        // ���üĴ�����������
    .i_acl_item_sel_regs                (10'b0                                  ),        // ������Ŀѡ��
    .i_acl_item_waddr_regs              (6'b0                                   ),        // ÿ����Ŀ���֧�ֱȶ�64�ֽ�
    .i_acl_item_din_regs                (8'h0                                   ),        // ��Ҫ�Ƚϵ��ֽ�����
    .i_acl_item_we_regs                 (1'b0                                   ),        // ����ʹ���ź�
    .i_acl_item_rslt_regs               (16'h0                                  ),        // ƥ��Ľ��ֵ
    .i_acl_item_complete_regs           (1'b0                                   ),        // �˿�ACL�����������ʹ���ź�
    /*---------------------------------------- ״̬����ϼĴ��� -------------------------------------------*/
    .o_port_diag_state                  (                                       ),        // �˿�״̬�Ĵ���
    .o_port_rx_ultrashort_frm           (                                       ),        // �˿ڽ��ճ���֡
    .o_port_rx_overlength_frm           (                                       ),        // �˿ڽ��ճ���֡
    .o_port_rx_crcerr_frm               (                                       ),        // �˿ڽ���CRC����֡
    .o_port_rx_loopback_frm_cnt         (                                       ),        // �˿ڽ��ջ���֡������ֵ
    .o_port_broadflow_drop_cnt          (                                       ),        // �˿ڹ㲥��������֡������ֵ
    .o_port_multiflow_drop_cnt          (                                       ),        // �˿��鲥��������֡������ֵ
    .o_port_rx_byte_cnt                 (                                       ),        // �˿ڽ����ֽڸ���������ֵ
    .o_port_rx_frame_cnt                (                                       )         // �˿ڽ���֡����������ֵ
);

endmodule