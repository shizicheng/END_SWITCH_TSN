//////////////////////////////////////////////////////////////////////////////////
// Company:         xxx
// Engineer:        yuqi
// 
// Create Date:     2023/07/01
// Design Name:     xxx
// Module Name:     xxx
// Project Name:    xxx
// Target Devices:  xxx
// Tool Versions:   VIVADO2017.4
// Description:     xxx
// 
// Dependencies:    xxx
// 
// Revision:     v0.1
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module Mux#(
    parameter       AXIS_DATA_WIDTH     =   'd8
)(
    input                                                  i_clk                    ,
    input                                                  i_rst                    ,
    // Eth_to_MUX
    input          wire    [AXIS_DATA_WIDTH - 1:0]         i_eth_send_data          ,//�����ź�  
    input          wire    [15:0]                          i_eth_send_user          ,//������Ϣ  
    input          wire    [(AXIS_DATA_WIDTH/8)-1:0]       i_eth_send_keep          ,//��������  
    input          wire                                    i_eth_send_last          ,//���ݽ����ź�
    input          wire                                    i_eth_send_valid         ,//������Ч�ź� 
    output         wire                                    o_eth_send_ready         ,//׼���ź�
    input          wire    [15:0]                          i_eth_send_type          ,//��������
    input          wire    [ 7:0]                          i_eth_smd                ,//SMD����
    input          wire                                    i_eth_smd_val            ,//SMD������Ч�ź�
    //verified_to_Mux        
    input          wire    [AXIS_DATA_WIDTH - 1:0]         i_verify_send_data       ,//�����ź�  
    input          wire    [15:0]                          i_verify_send_user       ,//������Ϣ  
    input          wire    [(AXIS_DATA_WIDTH/8)-1:0]       i_verify_send_keep       ,//��������  
    input          wire                                    i_verify_send_last       ,//���ݽ����ź�
    input          wire                                    i_verify_send_valid      ,//������Ч�ź� 
    output         wire                                    o_verify_send_ready      ,//׼���ź�
    input          wire    [ 7:0]                          i_verify_smd             ,//SMD����
    input          wire                                    i_verify_smd_val         ,//SMD������Ч�ź�
    
    input          wire                                    i_verify_succ            ,//��֤�ɹ��ź�
    input          wire                                    i_verify_succ_val        ,//��֤�ɹ���Ч�ź�
     //PMAC_to_Mux
    output         wire                                    o_pmac_rx_ready          ,//��ģ��׼������
    input          wire    [15:0]                          i_pmac_send_type         ,//��������
    input          wire    [AXIS_DATA_WIDTH-1 :0]          i_pmac_send_data         ,//����
    input          wire                                    i_pmac_send_last         ,//���ݽ����ź�
    input          wire                                    i_pmac_send_valid        ,//������Ч�ź�
    input          wire    [15:0]                          i_pmac_send_len          ,//���ݳ���
    input          wire    [ 7:0]                          i_pmac_smd               ,//SMD
    input          wire    [7:0]                           i_pmac_fra               ,//֡������
    input          wire                                    i_pmac_smd_vld           ,//SMD��Ч�ź�
    input          wire                                    i_pmac_fra_vld           ,//֡��������Ч�ź�
    input          wire                                    i_pmac_crc               ,//Ϊ1��Ϊcrc����Ϊmcrc��
    //EMAC_to_Mux
    output                                                 o_emac_rx_ready          ,//��֡ģ��׼�������ź�
    input                  [15:0]                          i_emac_send_type         ,//Э�����ͣ�����mac֡��ʽ��
    input                  [AXIS_DATA_WIDTH-1 :0]          i_emac_send_data         ,//�����ź�
    input                                                  i_emac_send_last         ,//���һ�������ź�
    input                                                  i_emac_send_valid        ,//������Ч�ź�
    input          wire                                    i_emac_smd_val           ,//SMD������Ч�ź�
    input          wire    [ 7:0]                          i_emac_smd               ,//SMD����
    input          wire    [15:0]                          i_emac_send_len          ,//���ݳ���

    //user
    // input                  [15:0]                          i_user_set               ,//�û�����(�ݶ����λΪ)
    // input                                                  i_user_set_val           ,//�û�������Ч�ź�
    //Mux_to_Mac
    input                                                  i_mac_rx_ready           ,//����֡׼������
    output         reg     [15:0]                          o_mac_send_type          ,//��������
    output         reg     [AXIS_DATA_WIDTH-1 :0]          o_mac_send_data          ,//����
    output         reg                                     o_mac_send_last          ,//���ݽ����ź�
    output         reg                                     o_mac_send_valid         ,//������Ч�ź�
    output         reg     [15:0]                          o_mac_send_len           ,//���ݳ���
    output         reg     [7:0]                           o_mac_smd                ,//SMD
    output         reg     [7:0]                           o_mac_fra                ,//֡������
    output         reg                                     o_mac_smd_vld            ,//SMD��Ч�ź�
    output         reg                                     o_mac_fra_vld            ,//֡��������Ч�ź�
    output         reg                                     o_mac_crc                 //Ϊ1��Ϊcrc����Ϊmcrc

 
);


/***************function**************/

/***************parameter*************/

/***************port******************/             

/***************mechine***************/

/***************reg*******************/

/***************wire******************/
reg       [1:0]     r_set;//ģʽ����
/***************component*************/

/***************assign****************/
//���
//assign          r_set                   =       i_user_set[15:14]    ;

assign          o_emac_rx_ready         =       i_mac_rx_ready       ;
assign          o_pmac_rx_ready         =       i_mac_rx_ready       ;
assign          o_verify_send_ready     =       i_mac_rx_ready       ;
assign          o_eth_send_ready        =       i_mac_rx_ready       ;

/***************always****************/

//�����жϵ�ǰ��ģʽ�Լ��Ƿ���֤�ɹ����Լ��ϲ�ģ���Ƿ����������жϽ�������
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin  
        o_mac_send_type     <= 'b0 ;
        o_mac_send_data     <= 'b0 ;
        o_mac_send_last     <= 'b0 ;
        o_mac_send_valid    <= 'b0 ;
        o_mac_crc           <= 'b0 ;
        o_mac_send_len      <= 'b0 ;
    end
    
    else begin
        case (r_set) 
            2'b00,2'b01:  begin                            //ȥ��i_mac_rx_ready��Ϊ�ж��������������ϲ���Լ������жϡ�
                    if (i_verify_succ_val&&i_verify_succ&&i_emac_send_valid) begin//Ĭ��״̬������֤�ɹ�,��emac�ڷ�������
                            o_mac_send_type     <= i_emac_send_type  ;
                            o_mac_send_data     <= i_emac_send_data  ;
                            o_mac_send_last     <= i_emac_send_last  ;
                            o_mac_send_valid    <= i_emac_send_valid ;
                            o_mac_send_len      <= i_emac_send_len   ;    
                            o_mac_crc           <= 'b1               ;
                     end
                     else if(i_verify_succ_val&&i_verify_succ&&i_pmac_send_valid) begin//Ĭ��״̬������֤�ɹ�,��pmac�ڷ�������
                            o_mac_send_type     <= i_pmac_send_type  ;                         
                            o_mac_send_data     <= i_pmac_send_data  ;
                            o_mac_send_last     <= i_pmac_send_last  ;
                            o_mac_send_valid    <= i_pmac_send_valid ;
                            o_mac_send_len      <= i_pmac_send_len   ;
                            o_mac_crc           <= i_pmac_crc        ;
                     end
                     else if(i_verify_succ_val&&i_verify_succ==0&&i_eth_send_valid) begin//Ĭ��״̬������֤ʧ��,תΪ��ͨģʽ
                            o_mac_send_type     <= i_eth_send_type  ;                         
                            o_mac_send_data     <= i_eth_send_data  ;
                            o_mac_send_last     <= i_eth_send_last  ;
                            o_mac_send_valid    <= i_eth_send_valid ;
                            o_mac_send_len      <= i_eth_send_user  ;
                            o_mac_crc           <= 'b1              ;
                     end
                     else if(i_verify_succ_val==0) begin//Ĭ��״̬����û����֤,��ȥ��֤
                            o_mac_send_type     <= 'b0                  ;                         
                            o_mac_send_data     <= i_verify_send_data   ;
                            o_mac_send_last     <= i_verify_send_last   ;
                            o_mac_send_valid    <= i_verify_send_valid  ;
                            o_mac_send_len      <= i_verify_send_user   ;
                            o_mac_crc           <= 'b1                  ;
                     end
                     else begin
                            o_mac_send_type     <= 'b0                  ;     //��ԭ���ı��ֱ��������                     
                            o_mac_send_data     <= 'b0                  ;
                            o_mac_send_last     <= 'b0                  ;
                            o_mac_send_valid    <= 'b0                  ;
                            o_mac_send_len      <= 'b0                  ; 
                            o_mac_crc           <= 'b0                  ;
                     end
                    end        
            2'b10:  begin
                    if (i_emac_send_valid) begin//QBU״̬��emac�ڷ�������
                            o_mac_send_type     <= i_emac_send_type  ;
                            o_mac_send_data     <= i_emac_send_data  ;
                            o_mac_send_last     <= i_emac_send_last  ;
                            o_mac_send_valid    <= i_emac_send_valid ;
                            o_mac_send_len      <= i_emac_send_len   ;
                            o_mac_crc           <= 'b1               ;
                     end
                     else if(i_pmac_send_valid) begin//QBU״̬��pmac�ڷ�������
                            o_mac_send_type     <= i_pmac_send_type  ;                         
                            o_mac_send_data     <= i_pmac_send_data  ;
                            o_mac_send_last     <= i_pmac_send_last  ;
                            o_mac_send_valid    <= i_pmac_send_valid ;
                            o_mac_send_len      <= i_pmac_send_len   ;
                            o_mac_crc           <= i_pmac_crc        ;
                     end
                     else begin
                            o_mac_send_type     <= 'b0              ; //��ԭ���ı��ֱ��������                         
                            o_mac_send_data     <= 'b0              ;
                            o_mac_send_last     <= 'b0              ;
                            o_mac_send_valid    <= 'b0              ;
                            o_mac_send_len      <= 'b0              ;
                            o_mac_crc           <= 'b0              ;
                     end
                
                    end
            2'b11:  begin
                    if(i_emac_send_valid) begin//��ͨ״̬
                            o_mac_send_type     <= i_emac_send_type  ;                         
                            o_mac_send_data     <= i_emac_send_data  ;
                            o_mac_send_last     <= i_emac_send_last  ;
                            o_mac_send_valid    <= i_emac_send_valid ;
                            o_mac_send_len      <= i_emac_send_len   ;
                            o_mac_crc           <= 'b1               ;
                     end
                     else begin
                            o_mac_send_type     <= 'b0              ;//��ԭ���ı��ֱ��������                         
                            o_mac_send_data     <= 'b0              ;
                            o_mac_send_last     <= 'b0              ;
                            o_mac_send_valid    <= 'b0              ;
                            o_mac_send_len      <= 'b0              ;
                            o_mac_crc           <= 'b0              ;
                     end
                    end
        default: begin
                            o_mac_send_type     <= o_mac_send_type  ;                         
                            o_mac_send_data     <= o_mac_send_data  ;
                            o_mac_send_last     <= o_mac_send_last  ;
                            o_mac_send_valid    <= o_mac_send_valid ;
                            o_mac_send_len      <= o_mac_send_len   ;
                            o_mac_crc           <= o_mac_crc        ;
                end
        endcase
    end
end


always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        r_set       <= 'b0  ;
    end
    else if (i_verify_succ & i_verify_succ_val) begin
        r_set       <= 'd0;//i_user_set[15:14];
    end
    else if (!i_verify_succ & i_verify_succ_val) begin
        r_set       <= 'b11;//i_user_set[15:14];
    end
    else begin
        r_set       <= r_set ;
    end
end


//��pmac���������Լ�֡��������Ч�򴫵�֡����������
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        o_mac_fra       <= 'b0  ;
        o_mac_fra_vld   <= 'b0  ;
    end
    else if (i_pmac_send_valid && i_pmac_fra_vld) begin
        o_mac_fra       <= i_pmac_fra;
        o_mac_fra_vld   <= i_pmac_fra_vld;
    end
    else begin
        o_mac_fra       <= 'b0  ;//��ԭ���ı��ֱ�������� 
        o_mac_fra_vld   <= 'b0  ;
    end
end



//SMD��ֵ�Լ���Ч�źţ��ж������ź����ڷ������ж�SMD����Ч�źš�
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        o_mac_smd     <= 'b0;
        o_mac_smd_vld <= 'b0;
    end
    else if(i_eth_smd_val && i_eth_send_valid) begin//��ͨģʽ����
        o_mac_smd     <= i_eth_smd;
        o_mac_smd_vld <= i_eth_smd_val;
    end
    else if(i_verify_smd_val&&i_verify_send_valid &&(r_set == 2'b00 || r_set == 2'b01) ) begin//��֤
        o_mac_smd     <= i_verify_smd;
        o_mac_smd_vld <= i_verify_smd_val;
    end
    else if(i_emac_smd_val&&i_emac_send_valid) begin//emac
        o_mac_smd     <= i_emac_smd;
        o_mac_smd_vld <= i_emac_smd_val;
    end
    else if(i_pmac_smd_vld&&i_pmac_send_valid) begin//pmac
        o_mac_smd     <= i_pmac_smd;
        o_mac_smd_vld <= i_pmac_smd_vld;
    end
    else begin
        o_mac_smd     <= 'b0 ;//��ԭ���ı��ֱ�������� 
        o_mac_smd_vld <= 'b0 ;
    end
end
/*
always @(posedge i_clk or posedge i_rst) begin
    if (i_rst) begin
        ver_val <= 'b0;
    end
    else if () begin
        ver_val <= 'b1;
    end
    else if() begin
        ver_val <= 'b0;
    end
    else begin
    	ver_val <= 'b0;
    end
end
*/


endmodule