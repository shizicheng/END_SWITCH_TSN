`include "synth_cmd_define.vh"

module  tx_mac_port_mng #(
    parameter                                                   PORT_NUM                =      4        ,                   // �������Ķ˿���
    parameter                                                   SEHEDUDATA_WIDTH        =      64       ,                   // ��Ϣ����METADATA����λ��
    parameter                                                   PORT_MNG_DATA_WIDTH     =      8        ,                   // Mac_port_mng ����λ��
    parameter                                                   PORT_FIFO_PRI_NUM       =      8        ,                   // ֧�ֶ˿����ȼ� FIFO ������
    parameter                                                   CROSS_DATA_WIDTH        =     PORT_MNG_DATA_WIDTH
)(
    input               wire                                    i_clk                               ,   // 250MHz
    input               wire                                    i_rst                               ,
    // ������ˮ�ߵ�����Ϣ����
    input               wire  [PORT_FIFO_PRI_NUM-1:0]           i_fifoc_empty                       ,    
    output              wire  [PORT_FIFO_PRI_NUM-1:0]           o_scheduing_rst                     ,
    output              wire                                    o_scheduing_rst_vld                 ,                 
    /*---------------------------------------- CROSS ���������� -------------------------------------------*/
    // ��������Ϣ 
    // pmacͨ������
    input           wire    [CROSS_DATA_WIDTH - 1:0]            i_pmac_tx_axis_data                 , 
    input           wire    [15:0]                              i_pmac_tx_axis_user                 , 
    input           wire    [(CROSS_DATA_WIDTH/8)-1:0]          i_pmac_tx_axis_keep                 , 
    input           wire                                        i_pmac_tx_axis_last                 , 
    input           wire                                        i_pmac_tx_axis_valid                , 
    input           wire    [15:0]                              i_pmac_ethertype                    , 
    output          wire                                        o_pmac_tx_axis_ready                , 
    // emacͨ������              
    input           wire    [CROSS_DATA_WIDTH - 1:0]            i_emac_tx_axis_data                 , 
    input           wire    [15:0]                              i_emac_tx_axis_user                 , 
    input           wire    [(CROSS_DATA_WIDTH/8)-1:0]          i_emac_tx_axis_keep                 , 
    input           wire                                        i_emac_tx_axis_last                 , 
    input           wire                                        i_emac_tx_axis_valid                , 
    input           wire    [15:0]                              i_emac_ethertype                    ,
    output          wire                                        o_emac_tx_axis_ready                ,
    /*------------------------------------------ TXMAC�Ĵ��� -------------------------------------------*/
    // ���ƼĴ���
    input              wire    [PORT_NUM-1:0]                   i_port_txmac_down_regs              ,  // �˿ڷ��ͷ���MAC�ر�ʹ��
    input              wire    [PORT_NUM-17:0]                  i_store_forward_enable_regs         ,  // �˿�ǿ�ƴ洢ת������ʹ��
    input              wire    [3:0]                            i_port_1g_interval_num_regs         ,  // �˿�ǧ��ģʽ����֡����ֽ�������ֵ
    input              wire    [3:0]                            i_port_100m_interval_num_regs       ,  // �˿�0����ģʽ����֡����ֽ�������ֵ
    // ״̬�Ĵ���
    output             wire    [15:0]                           o_port_tx_byte_cnt                  ,  // �˿ڷ����ֽ���
    output             wire    [15:0]                           o_port_tx_frame_cnt                 ,  // �˿ڷ���֡������
    // ���״̬�Ĵ���
    output             wire    [15:0]                           o_port_diag_state                   ,  // ���״̬

    /*------------------------------------------ QBU_TX�Ĵ��� -------------------------------------------*/
    output          wire    [7:0]                       o_frag_next_tx              ,
    output          wire                                o_tx_timeout                ,
    output          wire    [15:0]                      o_preempt_success_cnt       ,
    output          wire                                o_preempt_active            ,
    output          wire                                o_preemptable_frame         ,
    output          wire    [15:0]                      o_tx_frames_cnt             ,
    output          wire    [15:0]                      o_tx_fragment_cnt           ,
    output          wire                                o_tx_busy                   ,

    input           wire    [19:0]                      i_watchdog_timer            ,
    input           wire                                i_watchdog_timer_vld        ,
    input           wire    [ 7:0]                      i_min_frag_size             ,
    input           wire                                i_min_frag_size_vld         ,
    input           wire    [ 7:0]                      i_ipg_timer                 ,
    input           wire                                i_ipg_timer_vld             ,

    input           wire                                i_verify_enabled            ,
    input           wire                                i_start_verify              ,
    input           wire                                i_clear_verify              ,
    output 			wire 							    o_verify_succ 		        ,//��֤�ɹ��ź�-
    output 			wire 							    o_verify_succ_val 	        ,//��֤�ɹ���Ч�ź�-
    input           wire    [15:0]                      i_verify_timer		        ,//������֤����֮��ĵȴ�ʱ��
    input  			wire                                i_verify_timer_vld          ,
    output          wire    [15:0]                      o_err_verify_cnt            ,
    output          wire                                o_preempt_enable            , //qbu���ܼ���ɹ�

    /*----------------------------------------- Schedule�Ĵ��� ------------------------------------------*/
    input               wire   [7:0]                            i_idleSlope_q0             			,
    input               wire   [7:0]                            i_idleSlope_q1             			,
    input               wire   [7:0]                            i_idleSlope_q2             			,
    input               wire   [7:0]                            i_idleSlope_q3             			,
    input               wire   [7:0]                            i_idleSlope_q4             			,
    input               wire   [7:0]                            i_idleSlope_q5             			,
    input               wire   [7:0]                            i_idleSlope_q6             			,
    input               wire   [7:0]                            i_idleSlope_q7             			,
	input   			wire   [7:0]                            i_sendslope_q0             			,
    input               wire   [7:0]                            i_sendslope_q1             			,
    input               wire   [7:0]                            i_sendslope_q2             			,
    input               wire   [7:0]                            i_sendslope_q3             			,
    input               wire   [7:0]                            i_sendslope_q4             			,
    input               wire   [7:0]                            i_sendslope_q5             			,
    input               wire   [7:0]                            i_sendslope_q6             			,
    input               wire   [7:0]                            i_sendslope_q7             			,
	input   			wire                                    i_qav_en                 			,
	input   			wire   [15:0]                           i_lothreshold_q0             	    ,
    input               wire   [15:0]                           i_lothreshold_q1             		,
    input               wire   [15:0]                           i_lothreshold_q2             		,
    input               wire   [15:0]                           i_lothreshold_q3           			,
    input               wire   [15:0]                           i_lothreshold_q4           			,
    input               wire   [15:0]                           i_lothreshold_q5           			,
    input               wire   [15:0]                           i_lothreshold_q6           			,
    input               wire   [15:0]                           i_lothreshold_q7           			,
    input               wire   [15:0]                           i_hithreshold_q0           			,
    input               wire   [15:0]                           i_hithreshold_q1           			,
    input               wire   [15:0]                           i_hithreshold_q2           			,
    input               wire   [15:0]                           i_hithreshold_q3           			,
    input               wire   [15:0]                           i_hithreshold_q4           			,
    input               wire   [15:0]                           i_hithreshold_q5           			,
    input               wire   [15:0]                           i_hithreshold_q6           			,
    input               wire   [15:0]                           i_hithreshold_q7           			,
	input   			wire                                    i_config_vld             			,
						
	input   			wire   [79:0]                           i_Base_time              			, 
	input   			wire                                    i_ConfigChange           			,
	input   			wire   [PORT_FIFO_PRI_NUM-1:0]          i_ControlList            			,     
	input   			wire   [7:0]                            i_ControlList_len        			,    
	input   			wire                                    i_ControlList_vld        			,     
	input   			wire   [15:0]                           i_cycle_time             			,    
	input   			wire   [79:0]                           i_cycle_time_extension   			, 
	input   			wire                                    i_qbv_en                 			,       
			  		  
	input   			wire   [3:0]                            i_qos_sch                           ,
	input   			wire	                                i_qos_en                            ,   

    /*------------------------------------------ IP �˽ӿ���� -------------------------------------------*/
    //������ӿڲ�axi������
    output          wire    [CROSS_DATA_WIDTH - 1:0]            o_mac_axi_data                      ,
    output          wire    [(CROSS_DATA_WIDTH/8)-1:0]          o_mac_axi_data_keep                 ,
    output          wire                                        o_mac_axi_data_valid                ,
    output          wire    [15:0]                              o_mac_axi_data_user                 ,
    input           wire                                        i_mac_axi_data_ready                ,
    output          wire                                        o_mac_axi_data_last                 ,
    // ����ʱ���ʱ��� 
    output              wire                                    o_mac_time_irq                      , // ��ʱ����ж��ź�
    output              wire  [7:0]                             o_mac_frame_seq                     , // ֡���к�
    output              wire  [7:0]                             o_timestamp_addr                      // ��ʱ����洢�� RAM ��ַ
);

wire                                    w_mac_tx_axis_valid                 ; 
wire                                    w_mac_tx_axis_last                  ;
wire    [15:0]                          w_mac_tx_axis_user                  ;
wire    [CROSS_DATA_WIDTH - 1:0]        w_mac_tx_axis_data                  ;
wire    [(CROSS_DATA_WIDTH/8)-1:0]      w_mac_tx_axis_keep                  ;


assign o_mac_axi_data_valid                = w_mac_tx_axis_valid;
assign o_mac_axi_data_last                 = w_mac_tx_axis_last;
assign o_mac_axi_data_user                 = w_mac_tx_axis_user;
assign o_mac_axi_data                      = w_mac_tx_axis_data;
assign o_mac_axi_data_keep                 = w_mac_tx_axis_keep;

/*---------------- ���Ȳ���ˮ�� ------------------------*/
Scheduling_top #(
    .PORT_FIFO_PRI_NUM       ( PORT_FIFO_PRI_NUM )     // ֧�ֶ˿����ȼ� FIFO ������
) Scheduling_top_inst (  
    .i_clk                   ( i_clk                )    , // 250MHz
    .i_rst                   ( i_rst                )    ,

    // �Ĵ������ýӿ�
    //.i_refresh_list_pulse    (  )            ,
    //.i_switch_err_cnt_clr    (  )            ,
    //.i_switch_err_cnt_stat   (  )            ,
    //.i_Sch_reg_bus_we        (  )            ,
    //.i_Sch_reg_bus_we_addr   (  )            ,
    //.i_Sch_reg_bus_we_din    (  )            ,
    //.i_Sch_reg_bus_we_din_v  (  )            ,
    //.i_Sch_reg_bus_rd        (  )            ,
    //.i_Sch_reg_bus_rd_addr   (  )            ,
    //.o_Sch_reg_bus_we_dout   (  )            ,
    //.o_Sch_reg_bus_we_dout_v (  )            ,

    /*----------------------------------------- Schedule�Ĵ��� ------------------------------------------*/
    .i_idleSlope_q0         (i_idleSlope_q0)				 			,
    .i_idleSlope_q1         (i_idleSlope_q1)				 			,
    .i_idleSlope_q2         (i_idleSlope_q2)				 			,
    .i_idleSlope_q3         (i_idleSlope_q3)				 			,
    .i_idleSlope_q4         (i_idleSlope_q4)				 			,
    .i_idleSlope_q5         (i_idleSlope_q5)				 			,
    .i_idleSlope_q6         (i_idleSlope_q6)				 			,
    .i_idleSlope_q7         (i_idleSlope_q7)				 			,
    .i_sendslope_q0         (i_sendslope_q0)				 			,
    .i_sendslope_q1         (i_sendslope_q1)				 			,
    .i_sendslope_q2         (i_sendslope_q2)				 			,
    .i_sendslope_q3         (i_sendslope_q3)				 			,
    .i_sendslope_q4         (i_sendslope_q4)				 			,
    .i_sendslope_q5         (i_sendslope_q5)				 			,
    .i_sendslope_q6         (i_sendslope_q6)				 			,
    .i_sendslope_q7         (i_sendslope_q7)				 			,
    .i_hithreshold_q0       (i_hithreshold_q0)				 			,
    .i_hithreshold_q1       (i_hithreshold_q1)				 			,
    .i_hithreshold_q2       (i_hithreshold_q2)				 			,
    .i_hithreshold_q3       (i_hithreshold_q3)				 			,
    .i_hithreshold_q4       (i_hithreshold_q4)				 			,
    .i_hithreshold_q5       (i_hithreshold_q5)				 			,
    .i_hithreshold_q6       (i_hithreshold_q6)				 			,
    .i_hithreshold_q7       (i_hithreshold_q7)				 			,
    .i_lothreshold_q0       (i_lothreshold_q0)				 			,
    .i_lothreshold_q1       (i_lothreshold_q1)				 			,
    .i_lothreshold_q2       (i_lothreshold_q2)				 			,
    .i_lothreshold_q3       (i_lothreshold_q3)				 			,
    .i_lothreshold_q4       (i_lothreshold_q4)				 			,
    .i_lothreshold_q5       (i_lothreshold_q5)				 			,
    .i_lothreshold_q6       (i_lothreshold_q6)				 			,
    .i_lothreshold_q7       (i_lothreshold_q7)				 			,
    .i_qav_en               (i_qav_en)				 			,
    .i_config_vld           (i_config_vld)				 			,
    .i_current_time         (80'h00)				 	    ,       
    .i_Base_time            (i_Base_time)				 			, 
    .i_ConfigChange         (i_ConfigChange)				 			,
    .i_ControlList          (i_ControlList)				 			,  
    .i_ControlList_len      (i_ControlList_len)				 			,  
    .i_ControlList_vld      (i_ControlList_vld)				 			,  
    .i_cycle_time           (i_cycle_time)				 			,  
    .i_cycle_time_extension (i_cycle_time_extension)				 			, 
    .i_qbv_en               (i_qbv_en)				 			,  
                                            
    .i_qos_sch              (i_qos_sch)				            ,
    .i_qos_en               (i_qos_en)				            , 

    /*------------------------------ ��CROSSBAR����ƽ�潻���ĵ�����Ϣ ------------------------------*/
    // ������ˮ�ߵ�����Ϣ����
    .i_fifoc_empty          (  i_fifoc_empty       )    , // ʵʱ���ö˿ڶ�Ӧ CROSSBAR ����ƽ�����ȼ� FIFO ��Ϣ 
    .o_scheduing_rst        (  o_scheduing_rst     )    , // �ö˿ڵ�����ˮ�߲����ĵ��Ƚ��
    .o_scheduing_rst_vld    (  o_scheduing_rst_vld )    , // �ö˿ڵ�����ˮ�߲����ĵ��Ƚ����Чλ
    // QBU ģ�鷵�ص��ź�  
    .i_mac_tx_axis_valid    ( w_mac_tx_axis_valid )    , // ���ڹ���ÿ�����ȼ����е�����ֵ
    .i_mac_tx_axis_last     ( w_mac_tx_axis_last  )    , // ������ last �źţ�����ʹ�ܵ�����ˮ�߼��� 
    .i_mac_tx_axis_user     ( w_mac_tx_axis_user  )     
);

/*---------------- TXMAC_PORT_MNG ������ ------------------------*/
qbu_send #(
    .AXIS_DATA_WIDTH                                ( CROSS_DATA_WIDTH               ),
    .QUEUE_NUM                                      ( 8                              )
) u_qbu_send ( 
    .i_clk                                          ( i_clk                          ),
    .i_rst                                          ( i_rst                          ),
    //pmacͨ������ 
    .i_pmac_tx_axis_data                            ( i_pmac_tx_axis_data           ), 
    .i_pmac_tx_axis_user                            ( i_pmac_tx_axis_user           ), 
    .i_pmac_tx_axis_keep                            ( i_pmac_tx_axis_keep           ), 
    .i_pmac_tx_axis_last                            ( i_pmac_tx_axis_last           ), 
    .i_pmac_tx_axis_valid                           ( i_pmac_tx_axis_valid          ), 
    .i_pmac_ethertype                               ( i_pmac_ethertype              ),
    .o_pmac_tx_axis_ready                           ( o_pmac_tx_axis_ready          ),
    //emacͨ������   
    .i_emac_tx_axis_data                            ( i_emac_tx_axis_data           ), 
    .i_emac_tx_axis_user                            ( i_emac_tx_axis_user           ), 
    .i_emac_tx_axis_keep                            ( i_emac_tx_axis_keep           ), 
    .i_emac_tx_axis_last                            ( i_emac_tx_axis_last           ), 
    .i_emac_tx_axis_valid                           ( i_emac_tx_axis_valid          ), 
    .i_emac_ethertype                               ( i_emac_ethertype              ),
    .o_emac_tx_axis_ready                           ( o_emac_tx_axis_ready          ),

    // .i_emac_channel_cfg         (8'b0010_1100               ),
    // .i_tx_mac_forward_info      (i_tx_mac_forward_info      ),
    // .i_tx_mac_forward_info_vld  (i_tx_mac_forward_info_vld  ),
 
    .i_qbu_verify_valid                             ( 1'b0              ),
    .i_qbu_response_valid                           ( 1'b1              ),


    // qbu��AXI�ӿ������PHYƽ̨�ӿ�                         
    .o_mac_axi_data                                 ( w_mac_tx_axis_data                 ),
    .o_mac_axi_data_keep                            ( w_mac_tx_axis_keep            ),
    .o_mac_axi_data_valid                           ( w_mac_tx_axis_valid           ),
    .o_mac_axi_data_user                            ( w_mac_tx_axis_user            ),
    .i_mac_axi_data_ready                           ( i_mac_axi_data_ready           ),
    .o_mac_axi_data_last                            ( w_mac_tx_axis_last            ),

    /*------------------------------------------ QBU_TX�Ĵ��� -------------------------------------------*/
    //qbu�Ĵ����ź�                      
    .o_frag_next_tx                                 ( o_frag_next_tx                 ),
    .o_tx_timeout                                   ( o_tx_timeout                   ),
    .o_preempt_success_cnt                          ( o_preempt_success_cnt          ),
    .o_preempt_active                               ( o_preempt_active               ),
    .o_preemptable_frame                            ( o_preemptable_frame            ),
    .o_tx_frames_cnt                                ( o_tx_frames_cnt                ),
    .o_tx_fragment_cnt                              ( o_tx_fragment_cnt              ),
    .o_tx_busy                                      ( o_tx_busy                      ),
    
    .i_watchdog_timer                               ( i_watchdog_timer               ),
    .i_watchdog_timer_vld                           ( i_watchdog_timer_vld           ),
    .i_min_frag_size                                ( i_min_frag_size                ),
    .i_min_frag_size_vld                            ( i_min_frag_size_vld            ),
    .i_ipg_timer                                    ( i_ipg_timer                    ),
    .i_ipg_timer_vld                                ( i_ipg_timer_vld                ),
                         
    .i_verify_enabled                               ( i_verify_enabled               ),
    .i_start_verify                                 ( i_start_verify                 ),
    .i_clear_verify                                 ( i_clear_verify                 ),
    .o_verify_succ                                  ( o_verify_succ                  ),
    .o_verify_succ_val                              ( o_verify_succ_val              ),
    .i_verify_timer                                 ( i_verify_timer                 ),
    .i_verify_timer_vld                             ( i_verify_timer_vld             ),
    .o_err_verify_cnt                               ( o_err_verify_cnt               ),
    .o_preempt_enable                               ( o_preempt_enable               ) 
);
/*
tx_mac_reg #(
    .PORT_NUM                                        ()      ,   // �������Ķ˿���
    .REG_ADDR_BUS_WIDTH                              ()      ,
    .REG_DATA_BUS_WIDTH                              ()      
)tx_mac_reg_inst (                       
    .i_clk                                           ()      ,   // 250MHz
    .i_rst                                           ()      ,
`ifdef CPU_MAC
    .o_port_txmac_down_regs_0                        ()   ,  // �˿ڷ��ͷ���MAC�ر�ʹ��
    .o_store_forward_enable_regs_0                   ()   ,  // �˿�ǿ�ƴ洢ת������ʹ��
    .o_port_1g_interval_num_regs_0                   ()   ,  // �˿�ǧ��ģʽ����֡����ֽ�������ֵ
    .o_port_100m_interval_num_regs_0                 ()   ,  // �˿�0����ģʽ����֡����ֽ�������ֵ
    .i_port_tx_byte_cnt_0                            ()   ,  // �˿ڷ����ֽ���
    .i_port_tx_frame_cnt_0                           ()   ,  // �˿ڷ���֡������
    .i_port_diag_state_0                             ()   ,  // ���״̬
`endif       
`ifdef MAC1      
    .o_port_txmac_down_regs_1                        () ,  // �˿ڷ��ͷ���MAC�ر�ʹ��
    .o_store_forward_enable_regs_1                   () ,  // �˿�ǿ�ƴ洢ת������ʹ��
    .o_port_1g_interval_num_regs_1                   () ,  // �˿�ǧ��ģʽ����֡����ֽ�������ֵ
    .o_port_100m_interval_num_regs_1                 () ,  // �˿�0����ģʽ����֡����ֽ�������ֵ
    .i_port_tx_byte_cnt_1                            () ,  // �˿ڷ����ֽ���
    .i_port_tx_frame_cnt_1                           () ,  // �˿ڷ���֡������
    .i_port_diag_state_1                             () ,  // ���״̬
`endif       
`ifdef MAC2      
    .o_port_txmac_down_regs_2                        () ,  // �˿ڷ��ͷ���MAC�ر�ʹ��
    .o_store_forward_enable_regs_2                   () ,  // �˿�ǿ�ƴ洢ת������ʹ��
    .o_port_1g_interval_num_regs_2                   () ,  // �˿�ǧ��ģʽ����֡����ֽ�������ֵ
    .o_port_100m_interval_num_regs_2                 () ,  // �˿�0����ģʽ����֡����ֽ�������ֵ
    .i_port_tx_byte_cnt_2                            () ,  // �˿ڷ����ֽ���
    .i_port_tx_frame_cnt_2                           () ,  // �˿ڷ���֡������
    .i_port_diag_state_2                             () ,  // ���״̬
`endif       
`ifdef MAC3      
    .o_port_txmac_down_regs_3                        () ,  // �˿ڷ��ͷ���MAC�ر�ʹ��
    .o_store_forward_enable_regs_3                   () ,  // �˿�ǿ�ƴ洢ת������ʹ��
    .o_port_1g_interval_num_regs_3                   () ,  // �˿�ǧ��ģʽ����֡����ֽ�������ֵ
    .o_port_100m_interval_num_regs_3                 () ,  // �˿�0����ģʽ����֡����ֽ�������ֵ
    .i_port_tx_byte_cnt_3                            () ,  // �˿ڷ����ֽ���
    .i_port_tx_frame_cnt_3                           () ,  // �˿ڷ���֡������
    .i_port_diag_state_3                             () ,  // ���״̬
`endif       
`ifdef MAC4      
    .o_port_txmac_down_regs_4                        () ,  // �˿ڷ��ͷ���MAC�ر�ʹ��
    .o_store_forward_enable_regs_4                   () ,  // �˿�ǿ�ƴ洢ת������ʹ��
    .o_port_1g_interval_num_regs_4                   () ,  // �˿�ǧ��ģʽ����֡����ֽ�������ֵ
    .o_port_100m_interval_num_regs_4                 () ,  // �˿�0����ģʽ����֡����ֽ�������ֵ
    .i_port_tx_byte_cnt_4                            () ,  // �˿ڷ����ֽ���
    .i_port_tx_frame_cnt_4                           () ,  // �˿ڷ���֡������
    .i_port_diag_state_4                             () ,  // ���״̬
`endif       
`ifdef MAC5      
    .o_port_txmac_down_regs_5                        () ,  // �˿ڷ��ͷ���MAC�ر�ʹ��
    .o_store_forward_enable_regs_5                   () ,  // �˿�ǿ�ƴ洢ת������ʹ��
    .o_port_1g_interval_num_regs_5                   () ,  // �˿�ǧ��ģʽ����֡����ֽ�������ֵ
    .o_port_100m_interval_num_regs_5                 () ,  // �˿�0����ģʽ����֡����ֽ�������ֵ
    .i_port_tx_byte_cnt_5                            () ,  // �˿ڷ����ֽ���
    .i_port_tx_frame_cnt_5                           () ,  // �˿ڷ���֡������
    .i_port_diag_state_5                             () ,  // ���״̬
`endif       
`ifdef MAC6      
    .o_port_txmac_down_regs_6                        () ,  // �˿ڷ��ͷ���MAC�ر�ʹ��
    .o_store_forward_enable_regs_6                   () ,  // �˿�ǿ�ƴ洢ת������ʹ��
    .o_port_1g_interval_num_regs_6                   () ,  // �˿�ǧ��ģʽ����֡����ֽ�������ֵ
    .o_port_100m_interval_num_regs_6                 () ,  // �˿�0����ģʽ����֡����ֽ�������ֵ
    .i_port_tx_byte_cnt_6                            () ,  // �˿ڷ����ֽ���
    .i_port_tx_frame_cnt_6                           () ,  // �˿ڷ���֡������
    .i_port_diag_state_6                             () ,  // ���״̬
`endif       
`ifdef MAC7      
    .o_port_txmac_down_regs_7                        () ,  // �˿ڷ��ͷ���MAC�ر�ʹ��
    .o_store_forward_enable_regs_7                   () ,  // �˿�ǿ�ƴ洢ת������ʹ��
    .o_port_1g_interval_num_regs_7                   () ,  // �˿�ǧ��ģʽ����֡����ֽ�������ֵ
    .o_port_100m_interval_num_regs_7                 () ,  // �˿�0����ģʽ����֡����ֽ�������ֵ
    .i_port_tx_byte_cnt_7                            () ,  // �˿ڷ����ֽ���
    .i_port_tx_frame_cnt_7                           () ,  // �˿ڷ���֡������
    .i_port_diag_state_7                             () ,  // ���״̬
`endif
    // �Ĵ��������ź�                     
    .i_refresh_list_pulse                            () , // ˢ�¼Ĵ����б�״̬�Ĵ����Ϳ��ƼĴ�����
    .i_switch_err_cnt_clr                            () , // ˢ�´��������
    .i_switch_err_cnt_stat                           () , // ˢ�´���״̬�Ĵ���
    // �Ĵ���д���ƽӿ�              
    .i_switch_reg_bus_we                             () , // �Ĵ���дʹ��
    .i_switch_reg_bus_we_addr                        () , // �Ĵ���д��ַ
    .i_switch_reg_bus_we_din                         () , // �Ĵ���д����
    .i_switch_reg_bus_we_din_v                       () , // �Ĵ���д����ʹ��
    // �Ĵ��������ƽӿ�              
    .i_switch_reg_bus_rd                             () , // �Ĵ�����ʹ��
    .i_switch_reg_bus_rd_addr                        () , // �Ĵ�������ַ
    .o_switch_reg_bus_rd_dout                        () , // �����Ĵ�������
    .o_switch_reg_bus_rd_dout_v                      ()  // ��������Чʹ��
);
*/
endmodule